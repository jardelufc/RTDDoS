`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YBwRMYhsWb3+uLO36i5qjZVrBTD4QC0vnrM3uSmnAHUNwfw7aJ6WZGMOfX/9IlXpCYBXeT0tQ5tZ
03BsJvkdvg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BOQeGLTF7erU9o/TklBDBKFeA3lfuvTdg25F5cUaa3nUs01it/tdgyY47L3GIKqsVfdIeFhT6EO2
fwTA3Jyd/Rj1IzSkUjaFUgaBR5SPloH1LSrpHT2DZhMq9yKZyMW2R3448wF1XoOtkj7WPN8JSAlj
d8tgVd0nFtED7Xrjlqc=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
B9eI/iNLJbhQ5nXVAgx7tK3nRDCZcbRp3KDbjhfa9xntxfJf+v3EL9pjGdRc9zulyldhLNtjbcKo
VBi9t6lQ1HaPFPa+XZNAm6BSqqkQ9qBooKcwVbaOCCHHQ/DJN6HO8l3BxEwdblvFzqbHeLvnyqlu
aXwakK5R/Kgn9LpL7J8=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
l4uqmKHhP0iK0pYIycYjRQtILbnmt/xorSEUr2M+WSts2snMZek6xATZKDox0a4VuL2ZEp52fQAo
Ny3gESpfNp5vXcY+DZiro/Yf+vMcfUqkzI7/ZJM1C9SkWjWUbU2gGrjpIRMs8PN4EHiozHS+zH6Z
1sIYcyoLXXdbs74zuPGRYW34dlOn9+ijdm9sgKrHjvLUsUTB/yq7sGUYU591FXBeUl1YOBRUQltH
1Zj+RAMFhmmtHKmdzkAMCXok7MQXz4lnZ9IE4+k5DnAmKXsPmB3nkMDUmasmbOPTX3zF8l9MOmcR
jOBgsjlBxDhiPWMKi/B2R6A/uUmEI2oeqKnkqg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O1faw3n0nSObaWIjyGMdbodhQlrYZt/mi9Nu95v5U6cB7VyxUC4tBLzy2IOZpQLJ57G4w1qhjIkw
QXlIfURWj/23bqXzDjoIijOjSHBJdKgOQHItonCyULa0I/iv0sXPBBEffA8ndvMFOWUkd3Cga5x0
ryzVRbBBdDODOYiAwpspO97YgfkkLQn5RhXNN4oo5okZPBxHOcoIPWMJteo3If3MBBrpKRFutcgB
nf8FTufrot8/MZhLIUVFTfHdycuKYdFrxfEzFzRobfHqvupopq0gBCnrGrVEQFE87ySeCMd2QNbc
bXpXNE+ItPeiNBKjMRpg2vMKjmroHXoaOcfsww==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lY2R6sjGciF0qz5EVR/Fh9BSbSDdGzAT0Fp8nbXR8cwrjyzGbobGeTAHfvr3KLCPhuvp71FuDg5s
25fPN4MmFfP09GO5TYxGObVYqCmCRveQ0ullgCTBIOUu3cvalnt9qWcqFLSQr45kZjp8M4C6TsQV
damkcbyLiSHi9tqldCNi5Y/NeuyIKcfri4/U89B7vBqLiU6lAlN/+rshTOsAAuANhkQJg89HlOxc
BeytQZ4V0wSAFW31hPMoTVA2AgQYkK44ofXgKU3l4sGfBv0PbUppyyS2a30WPNcK28Z+7Zx49ayE
+KiztG6fwIdq1ZYDH1WO8ShCdNUhutYl8ABwnA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 432720)
`protect data_block
5PxFusCvZp3vOAUZxnM1sIxqW4xT9StVtSU4Gq2KzG+Wpe95UcdqUovCv7AgSUWYOVu+t1E+EV/a
DZ06yZPfrsvV7dpncT9S4pCs8T0FQXAHDzov2spMSPay6SNzFVejKmFnE4kEToxfs16/zKDs8OOx
md2Clk6XLVFBq7fDmw7wM6J3lwUjH8N629ywJLWq8jGerS00emGv2jolSjjFLBMq7WgmAzK7+hyb
n/EO3meIqWJjimSjuEiIty5BlQtRFx3NrXGvp9Psg0gLP0hJpbciGFaSnb1DIyLffJJAqtIN8M07
sGL8YdVyT/jj75NmBW0GTs7BF/e5FJFZEr4j1xr4k63HmSqCUT6JNBGl/XkS89TwIuCgCiwbqe0j
1fZ9FR/qm4vBVsrHuLaqdzJfAlSxsWrRhqK5P0gImn2xZL6fmHTcVsuFJCOQWES0zYAJCytuzE8E
uf1DGKU9l9GwK1/f0MbEX92iSomL6UnIakv1zZL/NdqEf43/1lm8lmG+QOn59rczz6JpKPFZ1MST
eRiKZaf+Ys2NO6reIkvjV9+O50T3XJOS+OognuFbGNWNQxnCbdkysFNq4GDueLye6+BZ3xsVzJxk
oVXkuf4J67/DzbYkXJ3MTD3eGZRu1ih0Q9vqY5b/ul9v1zWaJc12NbivzEpHYuTJYgUy4964GJ9F
+ApwTRCWN+nIs2HTXLCChnUauSI6vtSATmBKDBsaUvsDdv/f1RmkRqCEspsecXyiyiDRJ7nOk1Y8
cUGx20stoU1GlKkYhyIPYkgJj0PCBcjJ79ww3g6tmUXA1WZnNCA7z9gyUONHS15Q7EBhDLPs9E0H
61s7lh1L8whX3EUlVwW+WQg8HmKYnPKcRcNaUhlfEYBmvlVwoCNwRuzgxy6RUv5/1i7VqxvCjNOP
1gZ0NqU95us8Z/XboX1y6rn9GQsasHJH0vFOaIZjBICyfMTTEKsB675BWUZizZilRqinPN22nZFQ
fUEx49LaovxsGUZUcAecxwR+2FjPSRHqvqAmcNDA1Vrm24Qeu7FWLUfjnihrISvhLv3Zo//0cofZ
qXXx4Vm4UTj6ZfITO6pCASMGGEW6eKY1Iq1fufc7Ns4SF5ctw6Klo1rhkQwrUztn2NNPeV4rBN7F
aBf3Lst1eTSMwYvZjgEYuxyfi6cM1+SXNxZ9YsmDKpRV9weesOvG0zxUyAJYHglqqtuJX+5kNuU2
5PixJKpTSw8WXbpRA/MHHINgvDI1ze6rgPyXA7lTPiCDBys9ktjSipwetkyy6KZ7XI20VZl5eWOa
VgdThaFH5WSW3quxJ2rkC3JcrRqUOkuGba5nyDrgLte6+AmI5OazFrZmTFnEnTH8KMz7Lj+ulRtH
u9EksgsMTKvh2CdXH0H2aLxhobUZFmS12RLWO0R383+ZpWED1/xTwybWCz+d+mVjIcUQf1wC/OaK
CsA1wf8TQqB2Ffqpf/IDDFKnowyJwlNVHkSKxGapmZO21i+96CJ+1/V8NHH62hT3yfMNGR4QTD7J
W7y1lx4b2V6Nb7JnMbX9bBAf1irFXq53ZldcAKRWei09tZjVBlM6CpItbNfuuucGaeopddvvRO+q
hYgLrFFRbb+RmZB+GeYrKuoM2BYc3zp/bboP5J57qDFyWTzvkFOpnYp3gYRgIvopGM2xfxYGElrZ
ffh/ka2JsDsidM/O1mqlcGc3+SeRoUuspzCxX5zRMJcbiywjy73xxbEgDqz4VhRTIq2HV5YY40z2
RWu6bCZUREPtbFAdoTl+cxLKx3m6rLBYF/YcVaV6zTwrQjLPtl/g2ad0cLs8gMt2fVkvw6hMvaYq
FwNnBQrWHzAz3krxxPDY4bPT5Vyq27lX85Fqd+1b7CQy6M6CbJ48PmyuygzUirKdPrNNZ3KadDag
7HeGXQzkqWsMRfJ7Fm+zx/1l/TPMkoJmgvyTmNG8H3rExWBsJWqDdKqRVzj9QUPoMizfhikkTxeC
Xyzy/1vSiZDf0FlZRRXsUMRICd7v0nhliWY/f8V3T7tupe16NIQUG0icUa+gGA1y3DsJuMHArM3V
B84pbCOj1m9da3JQ27/UqSxFBpZO6VsFGn1s8mnn2LfhiJygAIzrw9Xc/qiD8Zj8vHouHIkVWBN/
ttiszvuoC6Dx+9RGNvtaErFIw5wtpy2mOENiEMowEuR/Z8DmiLQpI8aabLGlPgzGZyehNDsbD+gc
hMHydg9Ddl2/y0Y1KNGBVgxE6I7UvS3lSvq8WG58iGlHpQxPrx0ZXOgVBCXPT+0COk/r8uAug15f
AslINLbQbWAeyzpB3tjWbty3OWVVj7utbWS3x75VJNiTVoIrZB6eY6rkAm+qOmm9o+Qbcqe/pSHz
HJyOnnVvlZDTIGLMw9AVc7t9yPOrZues8fQqaSkGQBzGAs1hI0FrN8KA7EZ5N4Q8VDwcizjurbL6
3bJuBPEh+1fCj3Ft5MeP62gRa+Fk/R5hG7tEwgc8N++NlBnKWTcWyjcibTwOHzkkh2GE45NlGDve
v5t+K60SQioN8Qc+TQJD8H6aliXRDjVRlC1SwLG//fVvRHZXITRVsuu7VCRU8QV4pWOI8QN0cXO1
ZkdaSBD2f0oOtP3BMnKvB9HHY6TYuOxWcxUn5LEFO3X3K8y/BHHypcKeZ6w11LzgZYYaDJ4Vp8rf
b2u6u4C7Q/pHc1v7nr8QdypAnYrBqBb01kymHsZhmZgROl5sttx827yczL6PE34Nd9IGn1+4ZYei
nH4u7M9DpWFcLA2LXuO5pP8L4fkjaqLBcBH8y+LKk7DV5lMuKTj1C7JaVkx7dNZy+p+X31eEb6t7
ZetMl4VMCF1BdIdcZt8+ATxTDVVn05GkWqAV+Y27vZOaIqZ+j9+bUhHYTnZ0bTSRi/qxcFg/f7iZ
hts6kI7AF1t6a9pAu+6QZ4kWm68Y2OQvh5nm/97Avr+VYhDR8rO1FmTpbZ3BSmud0/6lWrNVI2Uc
DKp/Waiy4J2pg9vuvRoQzvNOoXk5Vx+TfnrRFnd0FMV6LpX3nBsMXuQbc9zpSHT/yqPxX4bv5mSZ
liuyDRUKG6x5L3W+q5zMrfu6xLkzMJ0d29CyYz6w743rG3Zv3RUMIHM9oC0x4h/9/wAyuduLdZmT
dKfbH5FIks+yUcaoTnORm4E3ksjRke3UM31LdyK/N11JadQ5OTIh4y5IDGrRE5otV88/3i9eWNUi
fcLkE2fsIHH5hYPUVgt8lNGGYYu9m1yRMb+Rp8AjLl6EX5t1DppnEVXPsPSXH2kKnFKnZd5QM6lb
QMmwC+L1qPyQ2IpawbykUrDK2ksSYKUWXKAAt1nYW8DQzsEJUfi1j9o7ZxkflJEut2iem/yMAccq
IFxmCCliKs8I1rLBZCY7iu721IiwUpGAg0IpREI6Dq1JFpRlT8w2pzDrm6F2sl+LDwOmbBeErV//
xPlOpasjCOnBRn5laA49GgcJFyyuo/DJCRn/RvFKsnRUxU6Q52btCcQ+yNAhCLwsEaKCBalJksvF
hZasr3V+6EQZG96D8k9yxy/kBDEhJXrWF6SODI7//GbqEct31iAtCDWJtqZWSNS0LmPRNf8xyL8U
Az5VawgaQ5wjRy1eWFaUvcZYkBTUZLuaIPHr83XItb1ywxdd9CpyP1TzSnmcYaaONXKJfd3abzIX
T26xZN5yBeJEwt0Eczmh5zyLwfgovdfIqopJzho4iG7uA1zylc+4sYEbEuwCPjaurm3X/wdZm57h
6tj4xKVw04IigZ84AfLm90MqLVkU2Mq+tZessLnNBXkdtpmIJEoiKBm4aQ0KkM4CLdIVX7njigFp
h8XE6yFN6lUCvReN81efNgOIN7/cez8kaCJ20/PuwDZmuCYdHzWucknG99ZvgYoqHUlygm8xyCfT
0b7h+7HUQGnvp840Es/+vFofsvJaKCGnXUudzGowv2YXZMc3GDY44xabaFCLzfDA0vUHe6EqnKuC
TwgR2DRp+TGnAOB0V7kH0yRWWmAmzg9UJnzA86I6hkSuBudDEbrpTT2SmqQh/GxeqLNj7B74DKA7
xDazmPwJobsdff1ic/UwvlTerbLtxo+d+e7dxKrqJsSdJYSo3gni3bSl9Pc5kY3q+Dh+lkfJ35Ry
k5dFV/zwTGNMnwooOKm3WpZ0T/OLzRKrU+m9q7jxWJBZZ/Yct5CfJWyBAhi1Zh4o4NihKfVeyNDF
VW2lq9uPKwaq4iB0Y9G5zIQwu1uDPLmMfXsi0fhrNYIMYOZlOw0s6ovke51V1c1g5NQ330pPKp8F
KLaXB+Sur8x734Fv+BBe1wUWuobYsP2xGp2uOX5Ov8aHJvTv9oYoLJ44CG6YU77xLd5A5+2SpGch
HYn6m3RI2TFFdr4d11nbFuU7XQUJ1jC7xqrYhb1dnSNwqKqZXxcq6M0ESYFhQred5i71bdhYGVzA
5TqGnfiX31pb0+zrROk1FTkKUKZBDxTi7nChhcKp1otoUJgfm+ubMJ/t7zPayCvDsC19526At0HY
kcqg8xnlBn8HHNSyY5B/QeoTeQByRr1MwNR7k3lYf4fKinEDJcLTOPfAbdnZe6lIl646OtnxkSl+
IKtxUJBhQPY6VOt663zO1mZ6gG4fcNTxGyO2oxtt5Xvg/fRkr3h/ZfjT5s0jfCS2r+6LOTBu7I9x
wU7yGMchwo6r9fyCCJYV7Ha0qIjJ9747RtWv/x3U6Gu+fRpDGEbQ0wfkP2KUL7wD49ZS1z/4wh9s
16rqd9aVJLfcK+OudPIibqWBk4OVTUPEqeE342jAXF5clDOb2rY4J1svhRmlGKX2udTK0BQNVGY+
elDqxZBxw1CZFaa88ICnyYww1LBUlZEOcnlGeRR3th8tybRpHuf8r4zqzicbE5kqIDyqIMI3UEW9
5OmaJyb0ROj72XynFOJRcpt2pchbZWQ6GDOEnZIKCQEatY4iOyB7o0hNpiVzVnhEzz0aUMlrpNYE
JCt6HvQnbO09AgkWUQ/g40wOuOa6zgYz8+bqNKCwbYYCN9L/6qq6FQlcOpNds0U/9BCGc5AOWLFm
GXJPBVPQGuZSQRlidyEjlGvpdccWMc0RZyLGvhVXiMr+6Sw71bRgUIqjBwtmihKVB7+PH/cD8arE
2Xt1v3ecp/TymCzTg70NTRBw3pLG4fnB97DGdDC34i2BWaDbhz714qVnzGj5mm6H/HUePDmlXcpI
RNxkITsjnCB9qYS5hU6CBN0jTi3h8zfs9WRBjiA3lgvloHWx/lqPXf0iv1FTwruan4ffPaIETezi
Uz4MEUjqQLJsRDF21hOyn16cOKUl80tLe6jyglvzjwYzREIhacMHngf9XBSIkCIlWEqCd+3rrgLY
+R3LV43SxI1qeZy34z3vD92YAOsXPD+XfXpzlSYEDxoKu93PKE5jWVCGimTb0T+dFQvKRMo0ilve
ns6wWn1mDI9DjcxU2Z58h7Akp+pZRlCocolnsJK6pIkNW1CeYzSykM4xUz5DCxTT8STKW9BQGgDg
6RWzmeMuaHMJEAHwgMeGJVPFjHMU6QrF/fS29sJg0m8a7sqN8BJBuRy1zUtPGHorhKZbhvVeG8l4
Tl5BR0+J+0cmGVhplmkkivy1d4Yjkq1d53Moplu7Q0GQ230aHoC8HLU7RU0UZSHcqqO2QkpaN+1u
+scu1+kFfDv02VIjrw544LJNCCHwJNFp1Vhe9LNRsYzTJ7oUfR/u3pKRevx/e4KJS3i24QU1tcNu
IyTty2b90MzAS0NArWiT5qg14ZbVhdnfeCNATyS0Yuj/6D5J+/Uf50AeXqvWlmAsWa4P7AxxrMrx
E+APTKf8OkdUp8PVx/H5jVezqc4MWxvYH8TpZCWgD4e/8EJkK96Hwo5QQloNpJVf5qqN/oLPKUoW
/AwNHtd5Zv+z4SvcUpa1Ggeitq//tpmGnFazMVu0rd8V6V7mg3vu1SF6sZraanhGHLVD1ENsjjJi
U3zw2JvDxddTPI4RIjX6OcVivNsmXgbVOZeg1l1YT6tfXitjlUwHF33p1ox1OKIy4hJWnsBnv9J0
zpJ3l3Pp42WedpYO6Wu2f1vc87d2xFr4MiTBTeJe7c508/CqHgdwfT47pidUvJ61aUuPaycRBvE9
ZEUU5MSe3+AIxjoiAai1MFihrtRd+cDWF//O2zN5MoNKXnIejBxlpS90avznAlwzBvgFdtKPImyx
5lyqtesNguMWqNajxrNh+ySfqGzRI3FUo8EkF00OELHRPqodWP1bSEl4rRrMVeMFZyaC5qy5+OwM
LmDyGnwjQVMy76s8HDehzxmCMUrsqGB3SgCg/9LmEswADH/3QgikQoyEES/wXGItta5HdEG6ZKMS
BWmDjcvNE3YtZIroN1qyzUlnEtnRZAdBE1g1q/y6lqCGj8KZcUuW2s/wczwlzGWRrnM0W4Gefdra
KHlCAul9e4/zPomU/7wcVWPXZjDjIAUhY0ei7fjhT4jroSyIY5qsYQ83WigR0o74Oz5v09Pc0NG9
yLCboMtlWn3QR3vi8Wi5F+39PUKRkXTQyeKV9pH1JPA1r3WVIK9NPb4lhyVglUJcXJ8us5CT86uV
n7rvE6z1VIsfOXyyc8T4zty57p8YOpL3x1TV1Ko3W2QZ0wSIptfD8MUsJ5rC/QXk/4D/hh65TOoF
FqX2/nu/fCGQHvzOd3wmJ/tKXRSmTFNuySmD+AHQHzamFYOGsOiGytfScg7nqr9DIIjIN/KmFlne
QK0GVzyhlG5jeP5hRx6OJCCpJs8U4z7XT9iW89Z7az+yoH1mX0ydEhnlLjBZId8m0/ibt7RNsD5R
FffSDp4PQHS6bQE9z5lPaUVFMF5tsN9gy1t1e6atcepJAYTKCSmq+LsIcLsCClD5zUhUDPZlXvBq
gokNsgHmT8ckEJp4MRYTYPdT4nMcpeFOJLPjJyzPNa4xGzR0jQcuBPo7O8u1xH0V97yYSYjfzseE
eNFzqoxF385FHIaBbSe7my1Bjs6eZYrkPAOSYQmk88g1I+Ap5vNZda9q+gNUmjmVfsUZp+qQ6hxh
3Lc/XXG6hyd/pNIrKyIhLfGre/YWQIBBcAooCVY168FVvw9SykeFEPXIEGZlXNa9S+WFudfiKqnF
0OqhUEyo/YZo4DW2q6k6jfodsMNLeh+6W2T3pmwIXHjW+DShVDq4k+rRftli4kpR3BWunUzYjlL/
WbFr/Wz7k/txeyqCpophlmke4QJr6qsadBV3slhc2TUchuYmQrcc8A9YVQo6d6sVBjGPsi+NmebA
0WN8enVMPppdwhfCUSCDl25wP3c3Qhzbd2E4eS1gf6FFg8mahQ81ylo0iH3NpBomb3FKKDZAWrRN
xA0lxjmyBHk7jRCv+QURubhhJWjS/LmsuGB3ldoS5/Atvyrb2OlRUPADx8OxMV+Y+avG4hWoyEMd
jhtyHVX3T5+NV+2AlrQEv2RgZ5O776ryTG3f6JKV0WKm7hvMfXNFXJGYMZ19MEtiAbcuMGcuqBBJ
bHgNtdcnj09s8WnaqybwAOSRcjY5HYJYai/McR1FwPfAq304bp7cwIOIbz+eF5o4zfj02+ILcbvc
ACekUCvM/I/ZiQrqudI+7LDiAPbItgKlZCuhDpxEpn7EpbKRbLjgQVM1JYqa1k4Wguug571c3MMd
t/Nw51FrHcLg9JgxbdxijZZZzDwN0AQ+x6wONz9KYgb6jg+4PpkPiWUYhlLDgEz12uddFnvJQDW4
0E/xUitiwQ3exyXmTaAgIkGuydfTwWO0Ghz8ZNPwb0Q3VOuKfzXwanDGn/ncG7pQqORs34SK8fyf
KzUivs6IY0oITUEN+OGabwFBw7f2pQ3/VPvV+XOqJbEfxIldfurxbpn4BcDJ2r7CU4vWNHuFtPfq
WwNBz3Dvoof8Tz+N3ZVYP0UWYtV1Bq8xPYyq30wZz8089pQgwF/ggknYnfK7BEppOnEm5HbHbnPU
tV+C4xwUIEI4slZ1LmFpahBdLaqs3GGwl6XPmrSiEvMD/AJ23v88s0FBO9YU4Q/1NypmgDLp402T
VLwjq7p+Ro6UYWoc3tkPzt4OaAfqbO+8zFvYkdfD03IbJfDVCLEgr+s6bwfS9RuPcB/DXIeYCcBD
vL2WhVaAzXgPrBtgIdnSJXIvD67/KazEvaZ0KQDWxljd35ljXN+HqbV49QiBsM0YsYwtaV1R8/Ub
BIc7N2EyPSvrH28cwNhQgZe+CqLgqgRZGTHUZqxzoE4r+8pZ6ar/H3smGAi0+K7VNuiZhJdaGHvX
dSvoXPKtTvY28xbAbVSdItLRhp7B8O4KJ5i5CH5m/+knmDEGv1+VS7OIR4UCUgHV5pjnt+GT11QP
Ugqtq9eMZdFYqUpkF01x872pa3i/OfI/hGII/O7G2N4ZAHySZ76kcRQRHIYXCIfsIJOwccQO0b3f
3gAdrr0GYdn1Zjyui88F6VEr62udeWt1MAEhRt1hQLoSsmA6E23L0/4KyS9Zo62tTuN3by4W2D/b
/S58xxOvmQ/VaX/JuAHJxQChnpagRaIjST2a2fz2fbVq88pikYmPQtTAY+oXyzaMIoV0yMd/RaLI
GWTcxFW6iQ+PCyuCqpHJBXcnPw64WZCkANo7aD6DELDJBrXQbNMY6RqY6qcTS5R7biscZEk+mASU
A/rxtO0ZnX6TYqm3JrYBqyrDBoMze7E1uh5iiM/JBiDcue9PmM07fDR77AIEwlniPvkzpSgV34Fn
X552rJW7Fcxu3h9fnkBg4ovx0knZcfgbW3VbAAEUywcg/TO3IuYLepQQIwuyjAlGv5d1iPlGS4NK
qAXqfSR3B7G7Zioz6aC6O0kP1aAhYhm2HJ1pA+hRavTy0z6/LD2LkCH9Gh9RMSMqsj58jOfuUK9P
mwnZ75/2eCicsAI1PHZMlihSEzMfZdyQFh3hwDPDGsc1Kl+39V46iObut+pLPF+9AKTPQB7nfMz1
pqJW+Xkn1oj9bpxuMC+BIppriXTDa6bkaStwcDdRGGGAbMJ91wuHAuJ1vrJggg5bgmjjxt8R9HD2
E/qGMU2GOjop7QkohZRhZSI/ow5vlclQaqWhZbU8el+BkBAoUl2DR9w0OtzK6oPBfK2T+FhZw8AB
yLDkYwF4GJLOoy6SrDVrDl1QHBunR9IGZ6Qspi6vMCTUybThCcsiE4ZDRCjelVa4FuuLmYLGLhL3
GqT0v/b6J1C0ZWi2ITotg7uz0WaDje/AU3g87CD1bHlIIeHu7Iset1M7Tm3EYAjjqM1cwdBqonqO
XEACsrc0Dm3OKAkXC7maBwfDNtyzt60C1uwDXUlo75acVYX46233dcQRd/FjCb4/WSCRgtCDXT7W
Mvxn59dDuW2XpWxlt+++uh6PkqYXNuZQLAHGI0nrSN6BWhiCbILxvVGKP1uGGV0bjeyFbIqlqmjO
DbRT0dpUMuSm2naZOBfUcJ0ycEZA3K9Fm8oHwQZljZgPG4fIgo5i845smPGqU5Pi3aDZplUbsO/2
cbiuOiPLkDv6ACUZ46nFqqZv8LLVbSqq3zuWADu8575AHDnRXivSAcB4BXBpSCb45voA6NBAbQpg
jxvJAV456IrAD0Yr/awqk0pqlFYffjljDrEhJhnhG5BrKq9vOaFJqYtttPE5pReCwru6/mcrN4zw
JluN9VtqGzvibZQVNj51Csqajm3Hd7Kf+yF5RqaZZzPMb+vcELDHAnTCC3U27LuEQa0AbzE6z3WA
7wEm3A7/kfWOhFR7RDOHExUqhex71kK+fckbLgUjLlIf+zbsRJwh4aXXcNTrYiD0hMWs8+rNFyjA
7sCoy3E7u3fFuLDnak+d3Q72y1c6i2z1lqux/nWfo6eZsFxqvWKyVAyca6ZGAs/4eDJ4a+4HEz5f
HtSp0LCVmDzW7DPb1SLAErlOzCv8MQLNhQx9FP4Pl4eOx3Ucb7oQDD0TS+hmN31ORwPgja5Tlx5e
ZaPm7OrtovXJtX1oWW6wr56k81zd2/eFJhqSmXJ2QejOypSCamnQX6Y5VA3Vrz+51IktYqR3IoPR
UIOa23k27FwSOot+sQ5PfhhMyc8/eXiLwSiazOu4cAPJch9YjJBqG1lGwM48EkD8C9UiCGSG/Ykd
I64z0Y2DysnJpLjKt06WvM9yooF/q37hg8S80Hvuwhh9R6LRpXa5YgRUEbsjHEnApOhxlYVd1lU1
nCYfxtJx4I+QIQfnIBTynrSLTEkEK9L+fgRMGFTl2XdlbTCRbpk8VQEhceW53upcFerS0dhL25yx
LpaF6wxP3J3FDyP1s/zAhM4BUwPsi5uJ49IM7VTe8bLGQybZ0ln9KiriMOZ8P/L6vPfTEzIa5sFc
VRN0JtfqGb2wKrE0t/UISr2MLF2GdeLY+/O3Xc3VZxGiDp/Iz3bPIdy2oZS27x6wfgLe1u+1MgE8
cd7HXi7VdKQGdUyUr7Gfa/ija5yqVZF44b9UTXFFAhyQHtDLR6MK711a2wEzZTiCyk7FyjvcBjW+
SjF/OjTwiyAOhll77ndTtl/P5rPXpqnZgeSJ8DiTrY4b3fbrGnOT279u42Ytn1Ah6EByFhsIgHAL
gB7Res4hIGjy2r8n8feYVHbo7bVRryM87XZEzKeXPkfE2n/F7JGFxeIW5wP9Hx5K4flewRUwD6VJ
xShZ6wkBnRORUlP4FeCbTawQP5dEWsJpmZFp1EKqk22NFDOpP5VohDCKBHEOHcl2eMUZ4XOm6UlB
wzNT0FDECrzQ22LvI1e5BqHHH7XIt5DIDxiLqwBSu/5ffBy5lBGhAmRKbD+4KJXjlJ2xycC0SZX1
BgC5Q3B/mUiaku6ZypdPS+VwGwa/mFmugiAlKiXUWCqFrKhDFPLeikCZJNhaQW+eiA7XqByTRXvP
6CBo4Hny6WVybi046pP8HXSs33lsP4FomL2h9qqLB6OJfHpD1oL33htPjOudjZBoHO3H/aCWuWk3
QSxK4/fWX5/NSLjoiod3dOon74tIidVAJMUwv7HbB676Gxnn5OXjthV55SSnMxwgxvDtXzo7ZTZ+
mlPaC6L3wewsD34uJE9+nIPr7/nqGdkR+ZW+W+X7v6cUAAu7nY9fAwI0vHhTiwn1Iaj3r3lOi24r
1Cv3undu+mhQOkdY7d5HzIWglFR1ScrscIkIVNZRiiXKmb5odTsAXmgABqkxuJks+4VxrgEI6tbR
/KrSc6h1hCNfct6OcaTnkCpdn7D9oiFzubIKHh3ecYG98NcIKj0ykGSWd94fpnzYN5oaCliL5+8f
snZJwhPjmQW1IkDx8xqzNNtqqh1a33ia/8a2YY4LElJKBu557CSxkUFKAY6ss+ArKU4KrVVjAKCx
oQkzhyPkcjsLBcoc057YIDgmlZi1zKUaoO7453jIk1Um0FKW52aYeUyqbhB/S7Sxjj11zKwwDgm1
0t5y6Vo5RTAYFmDwu2ApLsGCzVSCHmgH0ykNQo0vEujMoazt5ULIIpqNugtHzIvgilUJP4OQA76V
5k7Ooa3NHQX2ddJ0gE/eEHpIhDFJYnS9VfJqfFMTPKHDJxaCxWRTyksguI9d7e7OBCfCcfovefqa
XHQ1PtCsBbIFeqvt4hEBoioVTtYoxRoMPzgcIRYcKRJbawlZtj6ol6U79x8u5DQNg971kIKDBE39
32aJj54njc1R3jQOU+TfcgqiGGQahW0zQiq4UtVb7LsjDNF8LgWD9E3cfkkU8Dys32OLg3+ra/Lr
TR/nResMqLNSHcVhNpRYDsXIT7Dn25P1JOl6D40PJzEZrm1mW6cN/vcnATUetdCz53FNugKqsLmd
pCgJL5PwOwluGWCBmKDepIn1Pu3yK76bQl7nS4z62BPHAKvo7FPDGVJEr/UudqbeQNqwmjyov/Tv
vks7nU4n6oni2ONz6Blg5iO2IZ2XK/QzN10y10vOkb5ZZTWsC0NWYaxlS9Ot0WrH6oiXrJSbx28E
IjhoTzcTZ1JThHTz2Ntjible8Bux7T74v7d11zvx1Z8i951zBTHOzWvPAeYVkCxdTnVsYEvXT1Ii
HDk8pAfav1BCHqQTk1VyfaS1QYS5L5W8DWMuUhqvZ6SlADGXnAIIWOTAtHavkiTXGNP7u7MMXUPo
Sqj2CJ2TXCGxnZp18GISM4fqV8vW59R9o6TD6mT4ft5xmZzw+uHEtaYdRHqqCehRZU9QAg2Eq3wI
7hLpdYioXxArgB/8ZQpVqBXCVrq0KZhbQ06gtsNf8Uu0BtlUGM9weZSleskvtpu5xkusbxTgiav6
99yhlb7nA9e15wV7fKaXCaIErh3j1a662NaiGuTWVVqugJCgqvUQn4vK0uiF1Dokl1+8sevwZ3dH
0/nms1HIbcYwgd4/hZ6d8y8vrzz6hKC5rkhnGCtBZPvpY3ZIm8VyerCf+uq8IvWf7X4RBWCpkpyR
HYj635HnbqliBgumuzRFD9kdzYRa8ZRikwnO7CWme0oiI9x8ix4v/rBBMRAV1cFrS5D+4r4FJw/U
7e4UqPbxFw4jWOv2AJqpComlswjhPYBXLTvTQElMZ4Hy/9bigCx+QAPjJbPTnQh18JbyJP8WGKKF
6rHfqwrQ/D7yRpW6FpvbC8+oDWnPeIEHR2ypCcBJ3C/LuKO4SC9EOWC9FAWeQ+rQxXrWugkh+Npb
S7LwftFjAaQqvhvp9jJD7Dqq7R+anYLjyIiDkZl922vOJfNiMZNsRt2+/HOdK5+IioVxZoZ4lJER
ZwZp0NVUjS6DStDY1lrn2SmBFUC4e0iqL5G3euuQvrJcM8kMuaf68B2cTR1pSv3Apm3EIQowgTBb
R1GvYe0xSocShkppYSSCGjiquSa9WTdyycO6gTiS3s56oW0Rgm4Tim8vA345NBc0Gj0LfFqe8X4J
9wZfDWPOHhr+Bet5ANc+8voRC8inWxfGmK9Pr9KqJ5l8n38zV6kYcDGIc7GDMSYE47XE8KdblNth
Of1s3QohEoHjTjuiQ2DCWWdSMYsFKs2XYabSPwGoBu2KXRv6QN297brRGoQEZixQQ4GbXlZvaVVo
mKRaWpJxccuJlyrKPHdkuavnbl9/qP23JUu0QRfT128U5B5vqSCSpiF8LiJLhvmX7B7CrNkrFLq/
i+6MDfRkBOwZdQMefzmeGKcuqJtjpblLYsSgJGDqxpjMkZk+s4NFrjpFQzg8Jx7qvvO/vtqtmUwK
lS+URn/svGtnwODXjQAMb6JtaxYQbsmSvjPGnPKuFEifoijptweXGhSXULDmql9jDXq29LDAXWoA
yTPCB2ayRdCpgtV/PSyf/HnUebbxwuDTN2NWI2VqEzYu9ro1KuResyziTnc4fmncYE0kLIZzG4V0
o+HQnCXkn2srkAWc2aEDyxP3gh3mkDpr9hYWjtQtmQXDrwtkO5gHbzTjPCBxYuzjcee/LfrI8bCP
b2cH+HskXZQ5C4u1wjQy2MW3ZVMKkB/pDb6nOq4S1bE8CAaBS+gCa09Mk0vspNVcV/l0lbISw1PQ
63xGsrZywhn7GVoKGQN/IxDgmcIdTv+yiQnt6mU5hvA1jqJe1GIT1hqDEOlzYYowYa9p+rZ4vpGj
sNKeByQvr76+3YPWe2Kq4dAzIlyKQg9ySL/r/Jt/REvESBuvrE9aET3RFHOtSqJoq0GrCeQCNrp/
UsSU062oG8ShaNYlvFO1g3KNL30cVsoP8ZdLpV+4LBs7+jo35EKOpaJZK9uj5ilxNg2DThbfgphR
fbkQKHKfgmJo67ZwOXiYtcYT2NVLRSjuZl3d8fBTcYyhfV78+Iwvc5bS3WaZJ2ywcgQwvvuzgczm
TmArCzrdWWT5L+OWikitR374ZK16KNE8gTIx6Rp10haMOvbIKu6uXOHsFHjC15bDrAgJueaTfOJ1
ydDT/dEQ25HwykIR1YtIGhWylWZMuIsLgpb0HzYhVFMUrFXKM2TtyNQI1pibOh5Fv0pnS3QsYTaR
OEHSMB/w5IrrWQaLlgFGDL6uKI9l1xsS5vSwvIljRusa48gSB5bJVDmywbUt5VpaXl6NLqclYtom
AgIPgkOB+tWfUNyUSSMWwEuXWfQmIOJ9le6g16skJNm0D2YJnOW5YRDFdovmUqrKXjozv5FSgS2r
UjmSUyKQ2JnJVO7vPoBPftDV5u6/ddWOQHT/01vrpQQNWW5xoSWqE2IzL5cAvc/e3ifQzVGijX0z
VciVZ5vs0DB0w20kHQ4n3OR8S3A9gzh8nlahO4opfsw7t8Q3mZk6KNDV9FwL6/1cHXcUDq0nEmmG
MOA4BFNixMjUUMUZGrtPvGGbo9tlCv90KfXD6DW8BVHfmbIRyNXNHumpcAQTZ3TDlB8xQuPvCKdx
dkHT5fB+CMq8O2zpQAXOCWMIgCt8eTkIVfGJJe7IR2PUg7wKi8zW//3+rGyOC2kUU8DCvFIUCuc4
G/0DaBS0YwOQYy+DvxW10wC8msK+L3sCybgcuF1ilaVyWTUDo2iLdZ/fvijncA19767bh+oxy/JI
hfK5h5n04Y9Q/MZlXGeKkSlqH2MuNk7ApDqaZ/LZFL2skjqh3onXsxXZ4lQB2oCriq5Er/lDiNRk
t6ApLjnDZsoQPQIxoQzUYv1SwNDpqkCiI1Lzc9tgilmr37Y3P2NVPV9waENe75cuXRnT5+E8T6I6
Ww5dvcM089poUeGSdYGRh/0g1yIWKhXvyg0RDO8KSyLVaAwDAjHmsgABsDMzl8KgE8GEGTV/MTek
m11CSVidmL0EeGaqr8LiksGPF1DCdeAM9X5m5Bejo02qvRU1kzqaHhZk9X6d90Ays3IY7xPNxtlf
xR8G/hl8p1YXOaSsXMQG50OD3n6FYHKRVguSrNAZ3hQtlo/8F0Z9EXk0rW0JZ8OTngjJAZTf0jjZ
KfaGXAJB2pKGUmsEYENqv5mL3kGPa8JeLRJGrwCfdVIkyxsQ3oLJxa+w16abiPqshbXI0r98pa7P
RK1Z9+lqsPHpDYG2W8ZEz06e243FtEENT3+EC6qBITuxZMPE3Ij7vumlHweumMxc/5Rvps08wUt4
cJEuFgwoCMU+pc2rtC4Pvh3XzyMbS6gq1VHbNGDkpwxLFli08diI8CZQ9uNTxYFwdQ/+oP/8m1TJ
JuWyB1svB5NjTY2AlXQeSSAp/ugnSqaZaQh83NSxqEZVJYw3jSXdO4w5E1kri6bRUUxMNB3TjgFL
mmAHNCSRWzGdSsL1wL4Khx8P2aeU3VFDVEh2qC8wKfMS50cQpgZMV+fxPeBmX3J5NiyiwRuHuQlp
b0uIsuI1ygJTThDHKAI6F+wc09C+vKFH+kxpqdhfFIP82XAoUftQxIEWHKaHJV4h/f6MM0cbgVpj
u+KC1YDunw/V0JxF/iNQK+Yx8TyHAQ4s4A83MQo9k+HcthGBpPRlJWshVl4wAAYMzdECHUx9+M20
NM4O+AqLpj3FWYGumZiI+s6PZQi2sPVGJEmJPcAKsnK7JxTb3LmI3wM8UQRUOm4UsUurcZpdldAV
TqcnHK/VHGoE7BfZkbea4NzecZbIMYK+ODRWLrRsXt/SIzn8czaEKmai0ifr09YjrAPR0S0Qb/vU
pQA0GSzTQenRADrrTAhkqVNoZO5tskEjOPoBWE2trsFg5MGm6pq1wtEJohZx3e5QBiGz5lCY+Xmo
N1i9xcM5CFd2oaykARdry6b+8mZf7z9bmIljndj+TmJww3bdshE53PxDewkAnuJtrCQ+3YWNUJo1
qcIE0NyPpCeu/NBYFbFvwUYsporFfpS1/WXgL934IRwVS16CkRDyTqDAYYK5TFkj4GBJ/A6CmPEk
odBGGWePPpy6E4ULxk+Zme167QAE+VPVa/9u+MsvaaEfZWBKFay6LaWKmJHiza/CjdwA4dJmaeX3
6ZZTuxPTFD5v3ZYdtrxImLBYQr/sLLKNGl99EfMey03qWx+kBojawXWwtvzJeg4D9GKT5FwECJR2
5j4ssu8zV4RGC9EtEk9R+2+4PE2Sn+V5v8IanEZCJJM5TJdDnu5phZRaSb8/pFSuwWUTqpSCsZ9f
lmRnoFVX1Xbn5nAXgDBFze3T3gnUBpClWWvdzYmhPAaTrmGt9m+5Z7HO5ZhRW58fm1zOR9ipqDK/
JPl/D0e/Ff6/Fnf/7OuW9ccMKi1kmOHy08OcxU+lJazW8kKbyP0xy8yH7VfWX3xSuCTPgoPRd2qW
Nf6CJUy8pVjNjo+G0SefBhVTIHqpCpc47GZJfVnX96qanP0dfHPk1nXYHoGscKKcs9yoWp1STn08
GESLJo4DN1sdhOg/g9e8Z4s3WndV+wUMOnmKnY9OmZ677AYjUg3DWVahPQh72qtNrqfYNgHWUyId
TcF+xAer+RYxu3MmluSbHBjfeA3hglDnnvQdzHbG4g7LVx26aY4bvJ8oPfNjVsus+Tl6VcxLjxit
/9+vkpA1r4XF6Szx8yklFOA8523c9KlBzdt+oxydwx9ChChlzmtjtgTtixFlzp3jWUK5eJgohCag
wOuyFdLp1MVvpxZhkHxsGmC4jZ6khdaHgaBdEKqwql9VC0vozps2oK5XpT7S39hdAJ5VfcM3oRE9
bg11xD1QdOw38XS3rfkYn3V0Dt8gADwMr7aajxTwnZEgbX5D6xCcnCHuPJNFGB+cBiLku4dTtRCv
jCB7nfum5Whxbsyi0oxgI0U4hd8zgMALdCRdDfWR5dggzMRGKf6v/sCHHTzVnjqesC4kgnMaEN2i
kNZNmYWWjaqhH4tSH6/cS78J+9YM2y4kEj/9c6EpNsFBS7fpc4+iCdjhhjYuFelwKKZzmEK7p1yW
6cu+hj6pT6kgt0Two2/TpbELP6at1gwqgXwTT8APHXdYwF55cXjxs+zev9GSDDF/JNAWjUBw04lO
Yw9MMsLiBvEF7zF3wULr/APaRhk8bNqHg6MZ8QuilH5hQYrRcOLTTNleHSd8HoGJRKIfqjMzefTq
aq4PQAM+sHRhZs0NUncRI7KXP4z9jX4srK1MV5frZghMaB2C7KdT4spKms4OUtvyqWZpaoQ7Bh6Z
W/QQ9LJ/MY5J0H29tz4BHDadEqAuR+l64fR2GthdWCFQ/02YJ95E0ugEG+ZJPSWTNnZggZI3/Rox
xXtcumyGTKxCgUSxCP6gy/Yorh1Ro0MrkB4UcZlzGrOHUAdcadbrWHseywGdFCuWllkxaE8JzNTr
Y6x5ELMvM/L6uQt2aD46UKIjX3D8Ku12qelJs6nHq2xAKHDuqrqqMM20q+t2UtkgSTKuSUpCXFF7
6723VxmK/dAI0K/G+fBKUAIrQTEUFULFUClSfv3SGH4ZYXPteJ90sBePOuUG5yeGm70n2DtNTOei
TGfnRpWxCIyp+C1rWj+zzUh88ed+BRdCS2Y0LheaoU1zjwy3HvzVuOC992gAMruTFE9ft6v6Qzb4
vhCMNq7n5xSCq4QlDf+AuFCz2g2a89N6GBqAOaitJA/5q6YUw72X8ULlweDoCfc50lFK/wJskgJz
Ig05qfn0gsYcPQqEqgw1C/ZkAo9pwdbkJh3sDsvY0twsOKldmEFCj7CRWuOeiearxBVJ1W9SL1jv
TPADnlfS7Qk6NL5FPSlt3P1tyZCVbxCQJ9h5ys/4UuJgECDB1hyeUlcDd+Hqe2hWQtIsnpPWhuR1
Ox5LZZBmOul79ILc/2gDNmpGh6YyuTGFEEd4752uNWgJ4rsla4Y6cGH/E8EFvzTlXvXn3/s0xkRd
Oj9xGLai5xlDBTX+7yto2QXNVCIxmUk9b4RehbPFrqHeti4dixF7FEMehOkSWLFkjVhS06cUgCSN
FNp9GNY1NLChkLyPeX7HBGaxWv4nCVfPWSbEqKiXDV88wcWBXkT3tQwW2PKJzK2JsyCuv+CHoITg
ZLzl2fV8I4+AT/12geQuLvfGEoptEBAmHTwZTuWutpnIt+Tc3VmoBoPWC1P6gS39Q0DKKIfccZp8
HD8LGbZC1d82duCgpKNf+p4XDJVSpiEc4ERMl2/1afv/BhGYuWZjnIocK3OmJAfNNYl2H4sOiymH
qT/NkbNkDlHjhEofUcizGGZAOVa1sloh3J+YBwx2DfnVqEOAVaMANviZAHIkeF90lVvYhenRy63I
vAN+Xe5dUUIdhO40SS+2URPJ3SN8V4vWEOXP7xB8Z+5r1LWSG23HdEX7FcQZtfiC0mvjRzdN8uyI
ZBfNCPRU8ixVfy4uFudlFeeh9A/gTsX3cpcfo2mGu9ZxRJMOiQHB7rgT12E38tQBLQj2G/7KBbxJ
plhFVB/1kKdzbL0IyTMI4ow/l3yRHs1+S5yWMKoDPi05baJ/apaJgBJnSmCcE2PKfhYIdwt2fdxY
nNF7pBTSWQWNtTyq/Uvq3JeCZXQ6tU9flhqLYvOcxSV2XH+p5sFA0AsVu4Z8Y7T9OweCoWKje+f2
Z7DnvQRpQs/qbtF/WXywhhwD9FrWE2abDY7GJqRpfUPIFfTnLNrh3UhbeEFHf5BkJ6Aw57WgNTWh
6ci+QywSJx//C0mGK9PLbBcR0t04Y3P2OT14quKpRXCqaYAlDJ9Wv5j6+qZsHaUMOntsDF/kaK5B
9cHMqLaLKxvZIXvMABQq2p0TQ00EBFFfLDJa5uuUDLJt4uA2FfJNLuNgVyQfibLksJyyy2btOXG2
pLPorEYevh181FYuFEWQLz+DGz+7MOdb9EeWwZsXkO9d3nHeiNbiFdIFBmSvXE3QVb8aj8zDl1kH
EtXgwWJOSMqOtNSoUzAqAspzCmr91ksSQlcLFxNqAlNKlEtDr/g8ja6L9toXz7KmIiAOMlIDIebj
qk5zsbK515OFsbIrWAFbAzPVbzxiTdTHcf77b7ByGMXHjCs8ZDn5Wt7rbtBmJIF01aPRMHfrmBU2
965ETPo2e0Kj+mqiCvtYeu//EaOTEJHU8Duwi/vnKvg8WxrayuxyltTfCcI6cwP7wIRA9JxU4chn
coIUzPbIWPSqRpSeKy/mmyhe9PlAyWuxg9Yu2Jdah2R/7jGy4xie/iO8f3ySweYdVmIWKr7z5wcI
6tR+FVyiE2vevH7iG2gICTOLxmER6uoBsqazgc64Y8qCn4DIAS0OlZ/4XYmytYkS4x3+TRSNWOHT
qEuQEZGEIZPSEgUQk83CD+uN1taC7GDdZTHZjTeBzKXl2NLdSAQTtglYEbQ9ZzsKEE6FyT244Fen
15rK+HvTmIuH00qFcw4WzALhyHY52eY7b64PtzWyaZaKzak/6/IRXv3s87VrBBv5YQP8OJxu7vmm
+7+n4YoBntA3Dszio4jE7M7/vrRZKIzv0AVT63OGIo6Z1Mrk5ePyNgHOoy08ZP5BXSYLOTKJf1qk
dRAGdUKYQ//cWOfix7aw/eA8x4haXqIesD9i4k4lEJccFPgb2SsQ8OI9nJKqUKYJwlMO9SSaCp2v
E5gHfGG0wPRpGOGU6NKo5UfV5TxdmN0qd8nhbJm54vLe2t6nlemKPdLlQgohb26bAyIuOpgzYgDX
Vmu5XY1iMIhTizd+6gh3yOGBqaTuHcpHzKhlQ8UU47h0OaCDPr5I6G0spTik/5o6zH9h99/jofHX
MoASU2pbIuRkKfAxc7zjVGDjivxzg0FfV1tnOW7Gg6TdxwsBlO232HGImTWme1X7DqB5dMBGj2ec
TVwhUQjjLUNU1vbjJI2Jrkh2fCkLHHDov5N6LEt1TOSllrMrnlaMD2uzFakMpmddrzUmASgM9aeD
xJkhgJHgvsZTWxPTU/eDbm6S4tN4PPQ5J6+vd9HTMuiOStqg+MAg94IuLSg/R6FQDE+/07xaAWkj
Voy4dzguaWwnw69Au2nQLE9Aqn1/hqcmTR/vbfW7DSHYW2PU265X966m75Qa5hBXzJPv1x5Zc3DO
omo1ZDAxuY+Xg40jMD5ErEWKnjjJTAGCg1dBFOZoUvkvNg44oIhCd+5MplfsKFCsK2NNlNmcDjEy
y3pD62mDADVzAhka7KDe3Wu7SWX3hQokZ6y/opFUt8pQfQwiwrE3Snmn95Sa9hAfAJel9z8mCSWg
9ItH5C0DFYclcDo0lrfOGE+zuUEzARoXk8DGQFy9XT0/zdD4KwqexQDn7sTtFe4f4gmrVwzq7dy+
C9foqWsdGRdfIVMTws6ZfAM5lwP4NerX9fITjxs7DFCme8EcUiPzYTxcVkmzyUkRhhxhNo2NIZQA
ddjo5gOj7sIwSJHlh/hAC5BfqeYesyt9jomyjSObbQKFtcFOIf21eODvicM0kFXkSiUHAzQ9Qz3f
kY8C0T6MrfikUrMbyrMMFc13nXFlKL7ZsZ9TB5NHRRuCLsdwL5HvGiKR3zHptmCBvWbBi4s5POCD
UGBuWpXdtmjEk0fudnD2mMrGfycnz9oLa+JsdwHNd6+fMa329xSMADrZoOdtkJiYse3Squvi7Y9e
dYAe7iPGHIuqxxv8qXdB5JLbyGMtAim6d1OBcrmwch3QvhBj/7tQ7MpxJ+Qmix/EcNQMlXc4w7LJ
ALZYEVhvjUEDmVZy8IdeCe/wMO1LWwZNlP92UdOmldAeFuQFrx5QV13YMeskOwHfpasUXBySZPdG
97bHIhccyXl2OghvwF+qFv9lJ+28or0NLKvwakxu9ULOr1IEZYNZ9BerJvQmvUa+oczNiPTEGEfr
DRRAHo8gqjCpxd4K+N8Emnn+8KZDcxgmBLFDxifxDtjzfELtj0TLO9g+VbAC6LkdNxjSjaQw90OG
WFIJ7qQ2tFzpoReGB2JvX+fULDWEzT7/XJk3cDbH9s4Pcb3JlT6CN7R/ZTOwm7/4hiqJhu4mr9an
XpVd9hW6SmMWeBGGbJFTDhONCFxCDxst3xhyscmK19QDF5Fbzl4vjT8R+uOiNN2MyJoUeMA9Ggga
H3EnyMlDKcNSs5UuEZDpKCOvXrBOdohtxywCByUfiBUPOLajMwR17WE7elekT5p/CWjeyJObhfDy
FDCbydkeyk+fftEgAXJmgEgkZKGdyJdoBANfG4Es1NWMxXXCvNKUXqvGsWBXrA5F03HklRvkmAzb
nnI8tv3M/BQazJMMUYBUX59G/vjkiqU3A7iNT9OechXtWeTl/66pUVlFqx/ioKA2eq/4tS1m69qd
gR3ahagx5UL6O54Sw/RbnatmmElK3crihmczJ0TD+ELvt0iNjifYYFfT9F/71WFAltB6M2Q/Es9A
jSfRR4aifx8UfauflGKdoR0h0d5eEnIJNmahXhLXkz5BS4jSmDIIfcTakDYOXaUCG3qSQbbQ6q7l
PPgvSil1hE8/p95TcUjctIZpE8qQSWCnCLbTLlO+g3tXKopmBGzYVFwDzbPjjgmJz2KYjy6hbpBy
mmO+dZg5RQ5dk6Bt64NS+9DS9+y3yuBZnFaPaujCAyTMBEDuyxU/Pq5ih4EdbHGm8meSXkhMCCUx
LwIStGfQ4dT8bWpKwS0IdbETD+kIt2DPdGCA1fcVj1/ScDTkFy6Rfb4yfRkAT7HIR5GBhyvzbkvt
4vzcqfAThCWTfh260gqbUDRqUFHZDajvIkQr/YPiO+aPtQKTjCQDqs9r4zXxzgChDosF64/UwDmI
u7AAFsI+tJylqNITPwPLEFRXGesslJmktDGnCZxMwrXYBS4V0wt3RdWc0oXZEJLUy/uhZ5cdBLUs
1XZD4kdtlQlRK9dP9+t+TrpmA/lPskd2sY+QfBywVzOiXXxGhnvYDQS53fcEaHrbLHaom9X6OhB5
C58Z9R/T1Q95gDklg57YVJsIS0TCioFSvLX9nXlEz1TmEuhAuF3jYk9RiVKyM4Jp4i515M8EmG+p
tcH0nMF0YqrsHDA+wkz78vINnEiFtEAbOvOEn1eExKsUsYaRzSi/9Qpeq4FG7F6i6JdKkvbE9iVG
1ltPQrHBJFhuxBsW+/UZ5RmgmUEK796/oQBckmCcJAdn39C/ywvgXJMuzL5SD4M6jlFeqomlXItq
Ny37P+Q9SXl6let5RIIqA0Pfdre7EAYqGMcTHLkDIPehwAjmImdgnQ2kXek2Mvi+YfQsdj8CYXvt
/FPMpNjZq+5XkjG4vkX2A0sN1qTNx1vplzdIewFqWN3TpesWxng6xbEV09aA8q7iEt7u//+akZ2s
L2X1MIdpKjsLcSqafHU9r87Y05NPJfKB19+pOLLHTRfsJ4b5FpCG5y+fx+H2Wcx/tFxcLn0r9ubM
k9cb8I9OHR/dPBczbV+frjtVbkTaXlrFURCF11XecnDN+Zw1nfb7FFBk2YchRfQUyWJD83ULYT54
IG5Vexk8cpX6hj2PpzGq4jbjreX0/NfiD7WHvGDq+uzYkruSFgOBsHR5hZTxWECISVQ4cI0IPRuV
NM7mr0EC1MWZkhVf6bHWMwCP4fv5lWpm/NFQaHoSrl7QRIiZ4Q2LOd98AB/XncIJkqLW5IFJG8gB
QZlPvREetrWaYA17A6ipdEazGIyBDZXTS+SCxBWCz7PRuMW26ywrvTrW8rAf/x2oXTvLLCYsbhoU
gBL9gR1oOJ07g9yKB8eIv3lqo3xd5amRIJEU4p4m1VARKFpSDgFw0B96EvIbz8Mvy/SIzzhDXfNE
Cr7IyQdt7C1KLnaUFZ05ZgLS6ktHCaCX4Em7+zdOMy4c5rwJhGiZ4jX+ei1KqWP0sKtLTM0Lz7AD
FK/j6at4xBz4NAyK+xWZFwc3Ko8EokWkrAAt2AKkPxIi0P1dpnV4PQsTkAOtnQwNPB/GsjZXMKcT
+iIDJkW1Ay0QkDKU8MVqUvWAo3PMLzuaJoD/z6YxVQkkBZii8XQxatGUsBzhE5zM/7w6CPaLedkC
A4qjmr1I54LG9pwbYu29MuEURVTpahUxsgztnLjVT2vnjAdqvAl7n9x4xNxVEtd0QvIk1ghNh7XZ
mWGF83RJjSSnsnCYzrSOZqNvGMbgFkX59q/58q1X3XdEC5Tf34r/uXDUsHw5UibaLUXI6WelXNU0
V2YyinN0fMLGxIieUZyWeh0qvdWpy4aztpJswLCsYtT6jUjQ20XbPu2SUByMy/tCT9e6B6S1uSD6
GGTF+ILhgWmG17IqsS4EtZowzAspHQPvz6togWTF0BMggxPhspmkFZymQ8m6DGJTeAlH7JVH+RKf
jxWXZd2evaeA5pus4GyUiwUcDI5FbF41/ES0Cry0ask/vOHf+oJHXKrkeQAQ6Qw4psaW26FYQYeo
ywzH/3r5MOJMbj8esBJ50DdJbXPSUvQiFMfVIR3vxs5mTOL6xpLm3xPxEV47k1JzAEOoctturEpR
jyhVRuG3GQGpQaVeVKxftvDqRc0DkrgRgv3ffEmjyKkfe1KxEdjDKgqCS54TOuYUQ2lNXwfkevIg
gadJ5nGebzaTYoACSt1u2G8Lsk2JKbmeESRJuII9PqEv45MW55cYWmAi875VTxA4u3/IsD5AEHe4
RPzlsC+u9t5bXMu4Wdv53fFP+y4gVPEp6tPR8enrPA3hekiTu7LTuLYKD4or9mIZS3N4ZK1rwLLY
k0pzh+wL1TDlT10mS5UO1ll2YSk49dX225aapCGXE8zTTn/jiLIDgoVOJ4v/TiDjpEfxnQSkYVMS
1Qw66ngEZYSXPngA9RON1aihV8TIaQv+mpc6vziWZ5OimSrGIdxEzq4MiYqL4OltmShxBRvE7ZSN
JLfEPsjuguq6ZrluAKpCSA+xJP+fpekvwh/2q9ssaC78dPALoh7d/pLzLXrGufVeFUxkH4LDf2KY
dUJhSSYuAVv8/8ipXmAMUMuFuS/unSD3CrEEN8kEXzu7OdnoqRTzdLmpHWbVdrQ+HKXcYIAPo7NY
p9zFHVX9tCBGh9EMRf7aC8plJjcJrGkXsFluhw/66JHiTDTrNBil5R/mxE8wPEH4eXl2bawY7MGP
Ba5mmlms0mwS0pGHUD5BLDqjCaUeeSZgZ9Up889Va7YGZ8LgdWtzWbBA1Oj4IzOXmr3FW1B8bdHr
rt4MxtCK883+pfCOJhd64FANJMF2293t2hpM6hrVbO1XmETBeYETk18cmbGwLmfKZqPrweUsJucT
F2qL36xsWb1nLJKME+cn1zet0Z+JsLuuTc6J1M9xjIUR2LEmuL3wqgCeQejPTH8wyAgMIdcFxRh6
mQrqUScCiiTNzoH5e+Vj1mgikmrxoQy5IkvFOWCYQgFsmG4SO9LD4oiijwQyFCihT186Sxugu1PW
2N70ZK4z1w5A2mVN9OKrzNciV0AbMTJCpwQqigjh7MwfQoElqi89KiWZnPwAQniMHtYMsHOVQB3T
JDkqmbOwrzcr0acKWzvGRaoommn6j7Uobrze4BASjyfb1nKyx8sF5fmAyC/MvwM19K1aepiQCNx8
XK5aT/jca3Si/EvIprcVV1aoP2+Omqod0fmRGzAU8tqwNmmDH2tPDaKa4m1hOzgZmPwgIsJEMVG2
Xq6cVhXVnXag9TBdXSsdrDvTx08KaQb//XJVwxwUSlL8cKq72eag+jNCahZnBjNG+ImeVi3kO4Wr
4P6w7FEeytZEZcuZDfILyTn00hUvZzZYpv4uHT256GCzteKx/bwxMHsfOlec9C0yCL4Frqc2Y6iT
qicz4VnRnUFO87ecTtOuzFdKVfa1MQGwjNaQi5ImX01f6lJiv6HBhWxEKGgK8c3IeKWyoCAQm5Ly
5WyiSdHMjrNgWgvh7GRQdQheVxsZeul4cHKhfWgKKlmXdsmaeWNoc+8vFmT9oPcBpZhPzLbaGlag
W396U08gJilwXPtxQOYgCqM5aidFePVDHC9TA949wDDUGdGUN4yFNAK7aW+AYUNHKztr3Uz2S13g
3iJQnwIyLaC4cwP7KcaGu/lUpK8p6tOQ+9qyT/0OwSRk/zTzJlOCKC3wPCKi53dZBYaxJQjRHE+f
1EKD4V23AG1AD9gSyFohW4tyX8clxMqY/UwHgboOmX+FZCeBeqxOcXK/djOB0nAAgmniDMTXLqqJ
Dq853mkSjyQUJ7Eyf5YxWynJiB+svhkbXA/RpYzRNGUTj4Y6vnSUnrKkn75FGsk4+7wDUGtYpq1j
2bZZRXdoEOpZh9efO9dfqwdLBSh2dX5nQhz893s9+8lOPbJhrpzNJ6QjGWJctefeNvZCl7q8N+q/
Z+mdZokmoWFCOtN2ao5IRQLTZPHaowK8YFym0EC903RMZoyZnTX9bwcvOz5wabNddyoU0AwmidMp
0YfU7wBEUJpfW9nB4ko3ECf9dgVARK51OSs/p7t6pGoi7guaJiaK/y1vB2OeHRpsujLkKGdduRJZ
kaUlovjF6i9iNX54Iyjo0Xg4ycgpsBTiUqfSYpRJhO036lrQ9DrkhCtr0CITTpkP5v2h6unOvkHH
MJ6yHuzo0tRF2otUgt9rXl8jRNHMLY2sMFFCc48xD5sQvkW33x9Tzn3/CVUAFjl9ojfHaLL8OJCO
goVI+UPuW2gQNZyHpimNZHw5AYXPMvdYTLVJIeIUiHU3hTNRs7+WrQdzYYIjDmq2cAx3tjEhDV/h
hEdArcO1M0p9BW1gOS5zuP2hRx5Ph3hd+kcrYEuksk+2/BwLTdYFMPL9UwqZBbRwjIFUw9fX0iei
gfKa8hZPz3gKqTHG2TAc+fjhDmH0JMAOYii07SxHTdA6qC6eXIjxSaSfEiZbzqaurtPd84tOs2/m
3AXia6xt7OEUyFawO8Zn5c2Xfzuda04JyA6nTAD+UfAkG3OFhDuMt6rkt4zyKJwCoE9GjunabAZa
E2H/CtWL08FjWL7yYQFXBD9W8sqob7MeBJzedIkrHBKbWvQBk15MT6+jBe1X+MrEkFozRwfDsEzU
yE31HD1LAbm2FTjG+STc5bOorosQ5+OKzkJI7ycPcn7XTY+Euqp1IUSJptfGMZFZDOrNGpYKPA49
tERAOZcteNnOaTPrvUj+72Yq8/fXrAtYcqbTqePpA2oIC56kQNmhojyLT2BejaQFezZUt3ANdpK3
n30dUHNJygeS2rb+zJvc2m4EL9iaKM0Ti4tEyjkwKZMaLt4CJdhw7/mD0MdQkKERLJ4owmrkwOrZ
xBiEPkqwaVxuBnRdwXSGINQhu/RrmZdknZf0oV4PWycpaWBq6dF8A06htNtOnaL2ynRmuBj9Kmm3
k7zgiPXZqsV4f9KdPIDWuWgrju75UzDjhMbygk6hNUmGPJCFqEcpXv8mHt4NSa/PZVtylkm4cpcq
SRV80NVkEKIqHnFS/0S72z9CdjyfbQJJF4N+VoyeC6BLLx0ID9x2tcx+XTuGRyuM7qTcqX1Da4sT
uexnQihUVZvo4OLfnQNBRsAIIMGhlZ3WYCNiuewK1yV6H17UiPq3r4pUVhGYbUhlEuHkfF4aQASN
TyxNHgvCo9TupU36tVguss9p4AkDsa3lb37Qudd9ma7K5LS5Rzg9kE2LOjUAo3iiyyZeEJC/OK1F
PB55i+Sf+WxoBKPs4Iy5fohrAhUJVZCIlPEUpvi3XlZ72emLZ6Rr7pQ4JcAWUrsLkngHLZBZHLU/
n8Er5zdLsee1ih5BoUBCnBsGA/b0gxuLV6g+3XNKcYAfqiMhxVxuX8gJFuz0SmMhoz2f/2bByceY
wUkc5sGj2ZPJHcyqg53I/u+kh7277OP5MOjXiH9IjpPhOBIH/7fZ5pll9i62mMBwun1cJPq7bmc3
fuqNbbc/msGI2DfBqA8v3lgIDbrrG1hiDifohVu2NwxIoHoufqqsAT/05cvUXodMruIqjmBY7vNq
BMVzc1FPYozxapR94hbLi/t7eHda+y35BZjU4g5zxjjheGrXkPBEVlvHOBsf0grZT7/eSQ+vdu9g
iV5MGAge5ZOe3s+qPtzFRAOjWi8kNwerdPZ6KUe+EL9a6JL0yZeAqAswcVlqCdNwSmPfJocGNtNP
iSUnUrv4x7OoXN9KXeb3EBMmjnH6nrz3CerwF+bb5tmAdYsIRKbL1OBysEq6LF5jJYuuBxytjITA
kLGJwZhIUgogP9rvbdGNv4p+VY6GXJv8zVxgo3nkvT4gy6QplZq7farYqoDYiSwZ9RMQEO7duOea
nuxl+lgFq3Sr6Rnm1hrWM28H+0XSPNXKj7RiEPIrFWaG1e0ym6k9Lg89LG/Uobiw1eJsA6wK4NZI
dLNbe8p9VGxU6FVDhJUZSxTU5jyiU7RPzJVVCcMuT4mnEeDvjCN6xb5MXqlw0PhQD5Uz/JX6RsWy
/0PF/So8N9Apvd0MaVsd7NkzyLK7/vbFueWo2wBx+R8/3iFl1RkR7KULIWAAWp9lI6JgimyxPAy6
SmzsRg+OhDdEGtYdbrJA0Nu6MTwRFom3sdHVbExuKv14NRnG1PvTSCh7KCyRH33B3/Mzy+oUt1jF
nEpwUGGVRRb7B90WXJ1GysVIP6IaOfGjerC5DaXWDQQTFNcqpE9HURDFxuO0WSRpe3i5oCaW+A7w
AkbcnGC2zYiqz77zRNh9LxKj4K+T5Ju81CmJ0KQIvFBW20LPoBULHjU3Yn0jztQvbzha/7xtM0uE
jDpZqAVZq9Saq7GCmT3fYTF/2ZcxcYRyUIz9gjvwJMUpqvINmV+w6er7ehM7KUeYPtOr1cqCGhGq
g0jXlTNFPePj5+ZDwRRx/tTN7tveoH/MUcqAnOs4sLSkxTS9GDDe5TjLHZ9HuOgpZNWS2yjvgTm+
gyhAvCZQxknyd3elKmSYoCWHsPiOQKADhJomgZ5t5H9RkltmUrbT3gHoAZ3GI3bC13h2FwMjtlk4
h+sJE8imLOFJJGCAE1wCw9G0ME9IDugJ1r7zCFRkcki+DO/7Uu5OHzzvzunSp2uUrOFwQZZQ5C4A
p+0av3mEYNieWiAymofeWvV0HcE83uB3zV46rtBL0hLndExYgGy5rjWQbwwzqxk2SJWIRTJQrypj
c63WuptHu+hwwK8SYzVYxiiDFn0TzlB4snu22zfyuoWJBM+XNRB8/GO1nFYUQeYxcvb2eavyzuiJ
+gj5J/MUwBi4i6pubr3wN9Z9k4PuLzmmuSBHmYl8LkMKDnTuCjLh4SXesF9C7+Kz/5YbBXrCmSWx
cpxe3vBUx+snkNwmyVWK4rR1nslVgQlbxJI5ZGJ19gSYMpfIywAf4TT7XP4CA1el2xRn/0HGsD+k
sZEnJn8s9Mnqv/1AmKKoi34S7j3wJWH8YgY/l/71XqEu3n5uKiDGR4GtTTsOfPr4b1FUfA5SX0hE
GsAh84WOrD5e0ZU7slTxSvm+kn4g/LSG5/xI0xH8kbs/MmwFZoHoyWeiLI/YLMSUqaLGiCiBNA9u
IqGn4IUJ5vXyCwX/rfrl3H+9Wk2C689SRWb2QGd49bOwJ4KZOpC667NroVBqMMR4ueSQlP7cu7d1
/W9MG2VFXffcLlFhpW8ut1UOaGI88Q7nh1wIq3XgBEQqf+ab+TbFBynwelDbi0i6qbT5k7MbDJ3X
drr5IBGYRHTp63fYOnpU5vAEJtZx1A48I16pk6gc4q7ABwyyyPayYzGfATLUrb6w/39syUVHuoLz
SsMwibiGiHYq6ogE5xpmA3LP6ySkxPHARxCA2D+8pjN4FKwXTTU6G5dfvv10HMKAhGpzCTPwRWUq
rxdKNwvN3Li07wDtaPPlQc0jzj4xTtfBmah8HHowXs4gdwOTjP/7iAMABu8CLrKvvDui0cCpk3e/
wFUCf8N3FbEcHsL0OuMnRu8nQX8blS0yRkgSJbpIxslyrMKMfIlDFxVhbeYsNWPvpCYH69j4UKaa
JcGQ20nh4jT7MRi0Wc1fPWBemZ5GSW9E1b0ZrQ9D50kceWmAUjt2KYRQnNWZIlIXpnWrsflva4i7
+u19ttmrtfOCs4ALnH3/OU4SqIDyFXYHg55NQ/5O1Fp4qKiCmpPii7t3G9/ULUgVuoKarQAC9LiP
Y3s8xr4Pn0QCacfKL7bak+2hm4R4933kIOUE3JlR76AJ9egLFSKrl5P19N66/SdX8YGARuYKQ7dk
SET3j5kG3ZOJxDVNI6ebbUToGHU5DedYJCkjd0KtHH1m3gahedQT6WGwqkg1cvo+EVBFttt1lz48
r0gDtAeSNMz4UCV/rB/7VF+3Khs20imo9zGVS6xY8f1Ey8SBDbKi3lu5DKH8eZ9CPBWpe5APxpT+
/XvHIP2D0QSHLAOVqTtuxLAsOV2T21F8Uk+bII+/7mJ/dq3fUiLM6U8Jt4qhAj0CHNExp7i2OlSB
Gg5K5Oh9X3+SCBs+2VwSZWrqz56Zz+yMC0XH++6t11BwrEQNP/7C0ZxqhlMK+AxcgpJ+swUWiNVj
YO26eNFrEflKmzxe7sjzKqpBPHfFswlleWiMfLDR9/fECcZphQ6nt/oAL/3bSMrJeTWRFQvtM/wY
lyEkaByH6uEI9ypJefM1dfxkMvmczdxTC8Evb+deVMAdfggmTocBhtnIjwJe2bpueuKAIKpcFCYB
dAJeuTLZEMLyrJgexi63dXOZiQer3aO8IgEIuKKqFzGSVHtmWJhueUN4JGlqpFRl3DIs0zQgtrUH
CEvfpEmDdwS9PX8EhMgTQfnpHe38W3LVtkbmcdu9oifbt3x88M6boxv0ZnTmPLzZjDJYWNc+qIvs
arSV3g/L+pWmwsSF/t7REyNgGLgbiSSmV2syfyNZgQgpMGgBJfRPjZihJvuRsmpmyJ3QZsRMYfva
+fu3svpisFUb+1Z7nBnpje260rHLv9LS86UMBFZM/xIsBMfz0KfS9q3ONuO3Y8jiHPBSEfKmjmc1
U5IYgxFARZCjnvctDJwTdOGM1V0FpNgCCBpvHTyPlGrXPD4oO7yTE4FDVk2YlkdzSJs+lU+4Lr4U
H93fu1gF7S/M9ig/QdAoncMytwaIsJNOZqtLcCF3+zZsheQGRJVi7ILpIcr2HP7yWO1J0kwMw/Ad
YLvBbBgHmk+8qYFWK8eR/aQfRujNw8uNgZaS8C63EEyNXOFVmyNTDUBC/nML2d/K/apBunzKv0aD
T+U/30arA227kYEuqtxKixAIdFyfHOV+ZEFCyiAERsG9jNfQ+iA0prZQ1SyeCrhRpHVVN7CGg+Vw
X3f8iIGWdkeLNvvFpvQu9dVyQxe6qIMIW0EO/0WOG2UofcnS35/pM3kn0kqTflR9X7LxZKpRJ0fw
5VoipCXifDw63bux+qWJYpCDrLeh8Pt2G3LTxmR2LGFBI/t7wdMZreOTPlO6836S6CGcHtXVa7Y9
fOdUuGjHSEbuD7tlahtn7YsLhnFSKZvuY9krfdrlLEqg1Y85DHIaOLgZ6GMuHVqk4Xi837vFqFr0
B4lnPlBJWfehjbmtaF4NW9yuOVV4bFgO+Er8aOTzLeu7FRlSs5cm+JjCN/0gURepNEOozBd63qTt
aiGNBBz+FEXnGDodOhsNXrCsc3F0QPW4+mx3cjm6JD1Iv+WsDroenu3cjj2Q50Z/qVgXmsKBGurw
dwynTm/18g6jgi0Fm3O0hnE0OyDSD5EVabDtc06WmqrvF327Wqec6LeyzXId+4XvNsdACq7dl7yE
iCSdPdHqWLBxmboQqfl1FvjWehOTmLMVhx3Yhz74wqC/T9hHmWSxHd42DrOFdT6pZLJsfGPxfyZG
WBu4eg2XmDRjHKugvlebTBD7Ju82Gx6dGnameU0LgCfkWI3sU5SGpmjnkjwc8VJXwI+lL4NpSCeS
OEt7R2B8Ieb9PlK+YXyI43mVarw+4de+sXtaMKv8njsneHdjXhJKRPcL2Wmt4dZshF4JvH+i4hpT
0IbB3Th8HOSAlOh4u/P8U5T0IschReAwXeogPGGrfd1FTvB/oryTqmUSc+lKTU3sWRTdag7CHdzF
eqTxK5SHDzooGgk33yy5halFQr27CdZW8T1lWHso5G5y9bf7yQgNU9COY/Al+JNFB8pixvT+dtix
0FChHz7UYtRHfYK4UNtluiA/JTTArAj1jmFTTajotdbDUoW3QA5b2IYT/YoEDlDB/kUZV15mlk3J
4k5w/0ROdkmFJltMNKOue9EablJfHrACamBABnB5kga+SWsnYqdrfqZBEEFrcuefshsQq2Ls1n7f
yWn4LqeYMkTHEfKxbbYF/eOFegWRP+UZh8yYSJq7fuOBKNBpKYGHxSz5JWei2R4JlDIaTPYjbD9H
+FvjTwl2AnyYG37bZ4T2YSOX7wIIXQQQS60WAIyA/TAzjtJnhHqCF7hcTCUjusj4ISa0ElLBIFKl
yzwBweacnk2fkMltuX7ENtDInZc34xHIaGb3OGlTWzf9mv6ZWkFZwN24E90rLeDP0n2xPhEflNZu
tEyTK4CYu40MOi0zfatv2PP9gp6bNXOAblPPx9/AYn/ygQe+zJBxo8FVWJXtTdqS4G+HjsKNI1xn
jZi2kUVqkZJoQI0zp2i3k0+UMGI5ary5yB7ufoBiUYYYx+swo2wdu2T1S64tg7wo/bA4yuiT/4gG
t9HJQePckElUPg0hqq7DavUwvBFjeMPZE3P4jDvTaw9Xlq548auVHVAX//KnHfIk4Vn8ijvxkplO
JfpnW2ds6XwSP70z6nEokR1erAq/RsxYBmHT6819+DjjrwTwo6j95e4GxJrkwwJ1t/qAIjq90HcJ
I+Y2QY95feusoS8qbNDtyTYQwLXqfixzOsaUCG8uWH6uYzs+sQkV5TZ3gVxY0HJIttXkAMPFbh8B
99hR2KkXc2C/vnXUSH2yZNlDzBRXC+xsrgWXGUMJ78UPNd86jHw9j2SNlOy7H25vTG7oJpni/pze
fURrsnhHnWeE8WvVyAokxClFhOFaf0AbtCPRo4cfdIPBYW3kStF8OKdA3fIJ6ZD+OMmoDBdH3k/K
+LrrK2s3Tlci6/5Jpdiy03ve3MfEo864E+lEnBhY+ymYNbQDBD3BoFZx4QYVQLlxIc2hnl9Hfxvv
SPZz/5ribgj9ihQxbnET7zsbowNBMVvEegRd+0uXM87npqbt6jVtpeu+/XsNOxteiaZWg5r5MrLr
l0nih9WM1hboWtIJN3SNBC3BjX1W9Xlaoodw16aYBkMZqSpIIwASAyNNQh5Q5COW5ELjAI6SbBSd
m1hVEOU9bXq3yayc03TZNcFxx/QSXO3I7hr+fAsngAY7YGwop+Y0CTUYm/IXg9hA472quBUuUMbY
YyBSr9L1DWPXMeSfSXxXNlHYcS21OexO1omgl9kgvJQmmY3dYCkAdBq+cOF1iSq7SLwOpbSycR9r
dzwD7tE5BiZWZf18CEP/wMddo1lxgg2Gd9saSL4n4eGV7WUtP5JOX3geFbPtYUB+940/6w93XfNk
2WhScSUncrVzIDAGiT4VaoRDjKXty4AVGph+AXAGhL9jweWxP/Ya3y63OBpkm7UTxmdcJktmC4te
G1A1vUxn7b8n4JV8LdYjrsfGhlc1tigTxjc5YEr85s/zGiyQhhTaAq+ehPa8R9HuJ00JTPbgCCV6
8bilfm/tCc0QR4mNx6q6Asr9rAn1tgV9ojrAy6oWqN5EaGjVGlnKEPWgybY/hB4VCJY25d+xblq9
MhEjUiYbaIOu4rPpiIpzeuUv+5+N8RkwtNRZYUnWGS18y7c0PuDpCAZPiEmUVtJtcGazcUd3cP6P
wJQJOJUAEeu4WkgnUilgSVThisWqUoBnukbo+Hbf3Poq32teF1UR/i8L4/D+AaGKO/ErKQLzMYEL
LDlYINF6IuHn5Zt+1Z322XEohkRMh35kJL4EgOLnNAeKEqD6anpeYNiVy9Q/AwqPXqsv747Glw2v
l8I7pysW1NKzmw+aftD9YHdW7dHZTYbd3xDlX4Q91cixkokcNariygd6zN3sNiBJLNM/c7SEuXY1
PybYWGgJIldhcihfSHAnDja5fr+xqv4URqtC0CEVEFlNpZbUeeXWvBsxmKT8VRzrLMukOGwsIkhe
s+YM4Ba9EMLGXYFzfqOamZ5+2CiuMa/14I3gEw9PGrR2GcHcwhDnOR2E+yjepGT4pWioJEKTLwoJ
o3/6AecTN7JCRBqntgS3fZJbLGoNbxgRQXmMrG+FYO/ve2Qk/0Pb24qLmDsHQRPO5SklsppphfdV
pXD2d9pczxxGXuevt3ndb9+vczeY27Pfx+LKegfd8nMT3vVxu88T48+WsA46Lm87xGRcZQxhbMmD
hAj/4qCSioG14S2XAIpfvHxvSnGuowhALHjajzKxx8lpc7wSCmrWDH3IAmj6YJY0r1JYUzaT7lD+
RW1gLjM7fGbEZ8+lzFcdeGkbHeg2fxoLc6Q9XMPWFNwGdvRSdeRHT4mey4xRMjUrtrqYnPlTyrOL
EENPA0tg806y3yWea8ZvxSh8OVRDoOvgBTw34WMWUgWmnMiGVj5LI6MbNCFUrb/GA/ZtX/YRjW3i
YaOGQFEvxLV1AsFFYT9nvUa1XClxIo6aKGTVG9TG84e23/MclRcnOv3T33i2F9S/ElOiZWOI8mOF
U4TVkcSpdQEXzqu2T84Y348rvokYODTl8AfUUPNDeJbuMl7RWaKOM/IqLFcwi5gw79kQ8gvz2ZHJ
77RyslCdSd+evJOByFmYSBZeGIDsS37q/hvWOqheR19P0B1Iw4CjrjUvaaGabzhHfXA5W+zhg0Zg
HrAeJ4RpOgDelQfJjgpvvcKoBhCXhprwTxF6S0vGJURS+WG/TYwAtqVObT38OqLYhJMQcXmzOuj3
klhC+OaKoEXvRQ1KHAMRYsD3nnnEXlgSVqBzXRMb4x862XsBE7kRwqDa5+GsObAOdpFL3T8mEWbV
w2C0by5v76U/+9oVvtdwPJh7Uq/Ju0OhBAV5eJ/hpWL/G28LFqznZZH42LbnUXNXb2vb90KfckB5
A6wPivmDV1HEDUzkKMDNj9cnSDqyfTVd3HibWKpMn+0wN1IhvRi8TqOv6a6YnkKXWup8tuRAULO3
xw+QDPIed7v5JaeAzZ2I1Px4+8weQ1lbxn3GmiG3kEd9SMgLhNaRR7JFNWMltlctEqIkit52zlsl
3ANExdiFpCJ4em7AN78NKP+LG6v8BrfzGOqWIHaAOHoqXUgoDVlIC7A5RfoJSLrl2AAHo2vsmUFh
QEJg7sS65M6At5jPhzCVyrvC0g75nqcG/6wXJCUqc7SKEZvgoE/Qu2y2vFpHZOHnD6Raf2ynHWu7
lFG4T6+3u+olcTUs9J+ZXWacUcnDD1CQZ5OQCXRA1A7PI0CU5aZiyGTxMfCQGPDUcqHJV08jspB+
KjVuegsLPOi/S4x61xoUzeAG0viawA8rLw4mgZCT86zKkyaeHWUxY9teDmNgkOK+GYoFil71GZ9G
gCxZkl4xs2Lebtp6WoNSxoS2vGIwU0SvoCS91AslMIQAYXac+MYwxeM5/eiCC9/2aXUSgYB01Nlh
MyTYrhpP8AkTj1YaY+puLXtdbmwX7CBUIoAZUdiks/PF15UyolVrGMNMPm7Kjl8885k4/bb82Ohs
7u3b4XunPSd9EFojAk9KE+VKb0UOd46QTBOtE7BZhJFBpqoorhJ/SNjBNqSKhSAd09P49YuXzcSM
QlNbatvE/+xCsqrygbLyJJzM6uJYSjE2tK0m33xZx/GZtsTNPxki/r7FP8IsbAEz7ApDNkMt6Jbe
FYIMM/G6SYc8/HTUm2yMXDCH7RdBiWPpUktiRqragi3XW0pZFC8GNtTIZkm+WbvRm0ko69OLa2iu
YLrv2PIHa+eSo9joMX7vF/+RySxAodt9PulO4O/Y/34FKudaTg1nnIXoNZ1fT2z41dnfujUCeI76
nk+GSpX+5muXkTVSj5gdAKVoSfBxMzJTXv2cZl1dJormxEde3p0lsRN5/EenABmoHye+fPoSQl1e
SvAnzxf2jP0lSflJ9Rs+I9XPWbLweZgMuG/MVCbAYnv2AQPd7ev2WFpcieosiiJh/ELGHTN5Q7yq
joGtC3RDnkWBuLWP5Fk3Nd3UN/qElcOyUcGp89Mdlbp1A2U/Inf1h9hbLa05x8wtKdXEIBY+kW49
O3/XIGImPHVb4JlfEiT4cInYQ9jpLPk/s0cOZB1uDFVdaopTN/QXZo2ONCTGr1xxL3QpEX/paU+2
FOP92ujojb7SSbU35FVC1wtfHESwQBjKHD6wPSaQkYjtzyQb4L2gxtJPAE1+qXG4d8iAeId8+k7i
tGEz8hai8kOVkUZglDbqtdB6+issXr4hSYxCKopI2jV2waSJSZMiSLFkjCn3E4roA6J5udIIFeZF
FIz3nwHTBNVeMDvbhCZO3PXDGTIFEoiUhqNm2ydEB/5EOENfKvdcMrjrFqcBUlgFA648rWRERhU9
coo1YIK4kyCxXxIFfsnHfMVB+Zi09+D3KwaXyAzCg7TNurd+bGgerdTceUV/AvuoLi+9PKdNNwHY
BuBVx8k1SLM+y1BFgZGc/O7ZiJr971/jtiCbboC5BlsPdudcQ7tmrmFjXSqIIpxLFJ0YFnALOsNP
s9MsbalgpTCLke8K58VliUfwifdEyOWroypIE0vn7kbIvxR8fcYLhcpubCGpRy+1hIcwkDNOqYLL
X65H5UV2wTpC/MmKgW40aGFJgfjXmtoKPl1vobewh9sy0doK88eWXJylTCAJjRsn6bU1OOY6JEWy
7EBKa7QI0tNxm9HesMR4k36nFHuk6IGKP56IJ+9LdCzQp2OE6ylwX74VQA8eEY+aoi1vbdYQe03J
s9l0la1A4I7mm6ljb53185Pgl2XJPM5mYbRn0VynwkUGMv6OwiBYy0ACnyVBnfsdz9lUJHe/DCAt
az/efL6oClPCTUGDUu2cwcXrn5wpF67KyHRYVqtw/KMSJtAjiW9rR/JxLCqjqI+u0SEI0ctVWvwM
tKB+ECOqFq1nfCk05osROOYe7NO1Aj1sw0VRzzTrQwrPJYxtK52+MuCw0+5dGyTEErnki9iNKkBg
MttZFTaeSMH4bVzTlxECfPNjI14cn+tHdr8a++ICCL3wI6Q0W2lvYgSlqobla70TPHj22+JUgbJy
LN2pRLWSBwwauQAEEfnEklVsiDiYRj+MwgRM5bXIygGhSZlVHGLDjehJ0vw2iPnLIjRwlviDZti6
IH8/MX3lreWbjk5oXF8TqS23MvoMOEBYTTVJUQpKRLqyXEFRraYIvBbVgpIBA3GDwXTp6LYc3HF3
m2Zi7Bm+Wi8TmjAywXpO0qYJD/coThEd6low8DWnBPLxuLjcW/cvtOIKqN0BzkzIIvzRcDreVYY7
ZKpeaWHPFWDcMVpgQT/bgEg9FymIMu+I4GpSRBzS8najLTsIl9/26hi6UxMhhb9SDTGNBwA0QeZ6
QFj2gqvHEhLu6Mdn/t1Y2/XnVqOyEM2zYzWRwdkJ4I+A6tRTUn9bOpicqoX9v8hRfl1Q99zzPy0z
KuKNRopGH2KlVPP+pPicce1HR0SjwPuxgh9pFpQjFy5fKZ1OqLG9kHzETSDM3A+IUzkt/cTnkXWj
3z2O/pS1MumnvmBpNgLxG55sL68xWWmXLAmvqkCM5VQaH4x0SdyEaMUiTHLTzTQLtzPt6ONWKRB4
JTOXka8xLHlkVUcXMjEGv2IRmrKHwuT9bFbw+ZQB5bKCpVXcbXulOev8u/ufeSWDDT2APtLk0C2E
Bk6cjfOEJe01PuFwgCs1XfZdrKhZx2DU6CTJ9ZnjCXxqw72Xr84j8k8H6so5OODFlPhHetJLipdk
ZtkrSeGGin6k93XtWksXB5p5APEgfQn+bqENv5RQIS0cYlLARvWJMAGp2dl1ECzQFI8zLcTPoyke
XYv2HoQF48rkGQC2lMRtkWgJutHMjbBz1kwg0PbMEky19UmK6yj89oUkHN3TTPootlF8YW3u/vWO
EgWVoPWdO1RJU8EKXQXVAp56crT7XtOA488303CK8RCAQmHDXqTC3G9eraCXmfHlfpI0IVlvgNRA
XYioV1TK2zpng3ogHY1ibpOTZY8GQVqlJH92FLc9V+tUW6ygZ2BxCnGPfqHNRUMArBvzCSNP8FPw
yJ8KASzio9P0H5OqIzwixesQRWXgaQV5vIZ4liczIo4IUtMWb1ZHAqbvGJ+6oLJ9xERIpYT5U/Bu
Iow+cJhIDQUrBN7pGWv84kAVzMjmofCIXtR8e20S130Fs3/QOk7NMShGYOKrPXpsE4OP0aPwQXx0
NlSZ9suRlAP9Ijn5FwRVtNv99il5s4lOmX5frxoX+MI/VTlARJKvwZfrT2AN5QH0MLHrge2HDiFA
6j+ukVQ0hWTDFY+DYt+R1CFp5inJSLqgnaJAsE56EruS8q0oWIUG9ieg4TJsqQWCridicUeMbb+6
oP1MF28hJ0Rg7WT6fZQJU5jz63kA1Bo8S0MsYqja7as4ueRrjiFHe6z56U4B1j4nabFuESIVXun0
10/hyHi2DONuBAD970tIlOAUM0AiI7DNRFzJcjsbF6ZmpsCrJPCdJNwEDGT9r6MBdo3ZZEnPfQqq
Y8vCT7mequulEY2MBV4ErHU8UyqrLpzri6Glm/I6KZ0PMkvG5FCxMTTmU1VinoPvw0qhp+4qVACw
Ti2crMZxfaHuyCRS0JIgy5935vi62d2NeLKNtkdL9RAMO7NsRQuX205f04aDj9Dqf3nookwmeSJ8
1akft/pSEPJtQp9YSq7davOc3xaWrxFKShyAfL2vuATFVkN9FoFPX9yrVRqQlLb6LSwgE0JWBC/D
aRFAf5s0KXO6mKAur3RAtM4UjfWRSA7Mw0WK/a5TBEi0leBUy9R8esVIr4vfiEN03u6YkwoJ1YlC
BONBn0hzdM87Pf474/u/oJQoLSv+Pgvd7NKnESpGxRK6EqMtgNU9oX0PXy5e3DphY36oggFC11Id
08PixBAZ6yj/jgWQslMWsXU/MDh0G2a1JBuK4vBE5rqrrdYF9FVpuzNgn4WIO6xlRnuSZ303xrzd
MatVhMe0hCRs4tf8P4BausNjJM8A2AWDdnbIMXXz85gtbyalRzruhEGuk9obzffQwSmqFFshBqZe
GiFRRwJ+IX3lMGNGYDMLiCVZGU6d36aYcLOO1myaIWWkrUNo2KtDgJOaI/N3sobJCzzLiMrorSjc
FBnny1X5XfSOdEcQwa83QslYj4JQW5NFzuYaFUL9eIP7E+HSuGZMOCmzr5l9uv+J3kUdHFhXJisO
hwYL9W8Wd3yBnfKZOvdNN5UGP6b0nsaXZ1kwcNu6rOn0OceEupXr3Z7yYisekDoKRA5hu7HElg72
FIye3/PI9TixF41XyEq9u8lFlpqB5bmrwKBnnduO0S/6rQourobDwkfrr4sAFOzgD3F+/oR/XoUE
idi+fXSA6W2glOmyB06zTwVet1V7R7QAjKq+7WFqh7RESwxW63QMuTX6fA5jmyxtIJnvFSFsE0o3
628HoCgwH9Ekur+9UmcuyJUIY0tY5RiXo93ADVIxg1OXaL3bv887HetvFeIlrPQDshPQEG9CvUVM
mRwJtQK6igTMtqQBcXL8fkm7Lva1YkWFJBwCKssY+IWKc4w0+CDihudJ7jRXtQneg7wU8ivTw9Jq
8xBk80y1EgVj23VWxvj2PLyqWtpsB39Y6clyioXEcOBKrbWE+70TMqojACMDQPTy27Q2OKutdiC9
atGi+LLs4he4iNhjvqq0KHZvOldjrW94zDz/GNxt2NJTe9Ya/VA5oUmjgFpjHXwCZncCJSxAxAnZ
zEY/Y8BMfzKFDZ5x/28X9uVryeQb530DvpcpHwLAAV3VcssnLuhGSmFgGsWoE3ke49PRByIzsmgE
/rNFTqc8DHbb2SUnEcmRpUew+82YtwaYbLgAUbN/vBAi6ZM0xP5Ky5j9eRl/njVlGfLMPtMXKQB6
Lua4acL6qwBq0ql2HZ3msRL7jfOpTeo/YyHsbhwTElZs6X1r7lVLoWnRXvI2Qe1iS7irp8iAh+fk
Gn5Alm2753gZC5N7nFTyAFVmmzJ5DEdlS8AV/ltn5JwHTSEm1Hyuc+jSm1iNx8L3v/5jau5hjDkv
hGV/VZT9ofxmCT7MXec9t6gsMaqG4DarWkRPbdUhcjXCgacdQWgjJx6ZcxCSqJt6mIYuFmzrEzaq
0xAm4J+RdzxYVfeLjJK3eUMfcU3U8cYyGhaH0W5SarIZeo3n7IAe2+ECcumXQMhMP04K7oaJ9Px5
y5Dz5RnGpkCD+KLRbxLgU7LTHgilVqpv7vpGNXeL5QhQPqgv3t/uEX/obs4r5KcZYylV5Vy6mpcV
74zlqrBEvxYEs7LQvBMBc3E+AZ8zcnwZ23xcx4e6UeHxkaL6HnPg5U7h1Rz6kuTbbRx+ZE+FqWSZ
Glio4h/J+XnCKXLmhINm9npniwHKmTBJRVNwBHnX7bY+9dA27rB2YUvvKFI7tbpQEA0sbeOQfiNT
ZeiZd8eKLp0BBxW1vdWjj7B/oK8NA5bwU23moG0ZThX9ANetguwCfun0K9Jux8J9EIOyO0VX0fM2
EDbRlA2Ii8E40CPH8Ir3aONlOx6c3MvQJQKSSbV6pNFS+S1qYXxe90DswDc/u9WX3SpTSX392Bx5
ewQRn/xJNtbBAv7OUhygQE7YSpMnqLRBCI8gg+rpnxms+IxwFshLLANYgacVhZYc54VE/1nyEb5r
HVpgzTF4UxfPcLe8k3Umf/c6ZR2pM9DdL5aTo8UB0GAjcRhJTQyhlzZiocmDI82iSkIvvsiwbKWM
Uc1hA9jdYd3jG2jdjdiIgdtTTZLdvS4/h0IRR98fQndxBP0HggyaUP1VXPKo4ZR+PWqH3gXZywlg
EojTBrdC+iNEB+2J1P0LWIZ+n2qPJaWATWgqV9rXPJee5riGtZW8nNNG5edYwWWYpc76vHgXsdMb
u3Jkay1NLmJzzRksf5DaSH2q1th6aWO11AQ18fosWicCsjScqqc9d2zh0G21PkZVguBop3tq1O6e
5dGtKmtIn/z8luU9wmFckUA/af2ZYH0N7i3zWbttzrC7G/cp0YZ2keZNseCTPPpVzMOmvMEUx/An
innnJEiXc/mgNARanWVNmlww63xkgj0+V9hIccu3mWq/dd5nsGdd5I7edLIicmQwCbre4Bz/pSUq
duNPgHSx0cDeVIzZ6MIpAVxEyJAsbBAHQiV075Er/bLk6qVuTgW4/QVBywtSjz+4P+93yH8PlcQZ
DK0Di7YDudt67jhfhL0cf00V2INlt2gxVn82upmmqHz0QBhzVOgm76ChIkoodxh8TukUsDyZOzk6
Rj8Lg64PjtxEEDmgN7CNQSD/gTRvGkpUoK3o2o3EgFwnfTFAapg7vyMydAV2Esy6Hiy/0U+2Rd2J
uxJWrmWq6UXLKk01C97s3dIT+tBOpniPsKaXWF3Z/vKo3YBkIRL4FTndR+ihLxI8HqvrVuWTlIFu
dldV2Qe0w7qZqOtc1NQQo/Dn4uRgNzdBkU/jyfsfwt/nACSXxTXnbHGlVfOh3lSVAQDZLtSHv7fr
hQYSntslLBfcMaBa9ZyQK9qruznatGubWI7M8jcSn5yfrdqApWEr+2ZFBRBaRwHc/osKUmskZFTw
2crYiKqyxhKSdlru9e3iE91UFOEA80HrPcnZSdTgaOD1LDzpQOFwNFV5xcByr23osBtJkoWLK00y
cE/EmMGKumP4yd6j9yQ76xJhNNoOHWKOFvKy0yWQH6IBzkYvKv1gT1ukpdHuxi1gclQ2H3Wr7WJf
a71jVT3tS4DWIdhGcEQkvrRcpl7XOjZqvkIZmpcgwJ5nFmpNlRj/7QfRLtwEJNTNxH7Qq0g5i5N5
Tfi5nVgrpw6WI9Td1Rw4uD9PSykMlLcJ4C1P3rL3+Ro9dJWq+GLXK+u2d8FV4fgmVxX12qrpnbpG
MJVluBDkfIaRJ2VnpakVOgcJGDytm/+5QeAbfswNaOxhDiwmzzE6bu9fzdfNJwxy3yIGdVsr/ENu
x0w8Fqid2RM3ptzcLsXpK3dCLyhUr4ePxS5Gx1FLbzXfP+Tj/oJ8ezcXPqVkiRVNBI6Uj0CN+UUN
IcdHYCnO2qeOLWINksCCvosyuwFlRgkTmPHmAduGVdBCt/fGTXEvy9fcjl9y+j7cHfjdErsKApa1
b83lqt8waYBQsDH4N9zI+g5sC/tpz/hya3BObQMcfgMKHKxj0QvuWVYvJjjHvHvRSMTAaUKEvb+H
BdzkDBvPHd3SZpBhiWKE6Uk2bvj8GLGRMVXS1idIvrqM/DFAV1JfoM4wQuUZt3hEAJAfyAWj2TgL
+Sq5qjYLtFQGfmSViYN6xeAknb4cqB+KLJ8u+aBRverkl9wQO6hVaib9YHnJJi1EyO7I2xApnSV5
g/Vd2BEghRoOcI6y3eVFd1XgiGOKqx7gIJ3K3SQ+z25O6JalkPa6+h4/1+5O6koWj3eoQUTTfp30
Bx/7oXTziL3RGwdTam9G+gXn+kfiMcZw1l7lJUej6MuWO7vw0sLZJB2flZbzMFPp+sZ8l9DUhjUU
0ymT3NwSZTzdF8jfB7+SBSQtdIIJrZE7gO4II6oob2MzctlvMVIKaU9hX9EJU5UAxSe/XbxU2K09
jiFTczCAnIn9BZ9A4n33fh7v83MbcyltObVAXMVYONQ7NXsDkwJFJbkVXDJ31lM7MEfQh5d0Cx24
VAgQLY+V9ed8/Sao2615fW96300EMYmd6gWrerTbgP8tMd3T1x3HZpdeJRIRv2KtbmXMucOBsi1B
Jn+IwMl0AtDuCQuiqW0kHg6e9mL1LiCfqSUXlP0VjLHp/0AvzzNouBjgjGNr2WSLYP0OKnVIUIvw
6+bR1gpxkmYddD3Xt8Nr2FKsArHhQxx3UcoZxKxA3KqmU3HVS9DoiLSCQ+TusfuhcwY0aGl89AU5
fK1TBd///2VKj+qYZP78lpD58q9tNCOWQnrLFWc4ENyy8uRXSkYwhrWK4KNaaWN9p2xJGpXkbCp1
rA1Ib4NA+ZRzeXM/XBHsAc13LxPJVqKvSucnVmnuDVa4+3gTQCAWZWPhJXkzTwECi6GEg1hIphFU
JHN79yloN3uzZdU1lxRUj5FVpfFtGC4W0ZCd/CVIxFtEbMxCRZHUYKyxx1mXG1KrsOh6cR6clW6b
KI2AHnIIOK1+2uX6dohD07otsAiebyMwZqheIYQF0t0m3MF9Zop89FTN5V1Y5YxCIyhN1zh3yk9M
dqWkHHczwSQRbrIXyvDZuxSJRPR0TO4cHwFJB+xYax0gpBDn+gEcY1s8WwPKRHStpaLJ1irOR2jI
jMPyJKH7WY3hY4n99bFgV/h2Lgzhp9lUfpbVLZftbuNZKpY9A6dyTw466K0cZIs5GDBUx6p5KBWW
gu/vpIUojfa9BamURiQmbvchP79jwNAhg8Ym1mtwn0rOOtGVmtND9s80LGe0F0qHPQAcTTytvfub
nxOpxeqyX6r8ly2QjCKfX63Y7WqltiFKbINeadslKt3Ba7eKttP+R0ScwHAtatt32AOsOdDhUYyQ
FlhCzOIRrbcb1GHoQbzbNhKr1EvWTco1x55VI47PyLkBnFkqqBoguZLHb3a4UC1OSSsGCMwn1OcB
WFOXgTV5ar0Lhpcho4B+7lFNaWVehXvFnAfwU19tg60Ocr609eVU3TvQzNUxqj46+Q3cLCXwJluC
Vur5G4tITlSoTPDpMxvO2z76J7rI8XfihemIlraLEIced/gAmVF63evvBp6lZkVyWdmYPEAgXlke
KDoZf5NGNlmkchEoI87iYUzT5vOZXo0mO0/1cUyfRPGva5bImXYCyQ2Iyoi/PxBqYU6mAL5gG6g6
7w3n3KY7f0S420ipiqxgcIdwODUxxCRmj3jZbzRvjFiSQJ1hbD/q1j3FUZAt2xjEYG7dHAwERlN4
mRrkG67n0LRHGrDdrOZRzULpVVXUhJQZARjAtBG2oUEnI2R6dc6phTZDaBrc+6sJ+vlSBk9mu9Vg
lUMVghvgtW7+xblP7p8jpcmsQqER8WShPkF8aVzkulC7QMBMAo9OG9iIQNPMmFXNFGpzoUiF2dP7
FNxo199mY3oBCKcltxTFnrwH1alPyaKJ5IZAL6qV/NlKe7tulXBszxfJ5XNpKRSrz0brxWN0cm44
onjZ+CXNtABLsNsf5H0eBLnVZNBcwpqOap+/lh9wbYxuBH3JdKyDMRH1KdSf9n8uEpctF7x6Ayds
ujHQ4uUdjyfEtS3/jrcktNgm/HULxLP/A7YT/VOe1FxyUBLnV5DudlVitXYpGPM/GgK1WeOV+nKE
b7laEcKyRIv4mwWjRaetpbdZ9Ab34nEn2CqBB9RBQALPng2/sFpOIpI/ORhDvU13CzWr0BF0cPZE
zP3zNP6j575ft+JhTZjQfG0NLi/8t3q68Mm3R9V2osq1vNex/GgTz+CnQiz6usT9F16UyDenLlT3
sc07dnfN1Zw9WXX/zHH1t15whU641+BmcBP/cxFScS6Xoytd1AgDmPrmmzj0IbQhi+DMrZAOcmkD
tx2AyMmUhu/ORpHwpBZfydQICeyQLWDoNdx3BtxKVn/rmQ/z8qbcnZFuClRtr1Avx9k7kYpA/PVI
hyjqfoRexn2gPml2FSHyv9ErMFTJx2+RsqsjHDx65GrLBgEFG4+E4e/QHeSnUnPtuLxQhWFiFw1L
lqftW+wbBM8O2aly92GmtgbFBEInC2t2W7f5aDvyYYHri/PsAs3b/HSI413Y6+/eOZjsld/sdT+5
a8xxNAuiwatgEvUC1nLOW4mlaUMN/BnW+9OAp9rjTJbRWYjip53mzWEEjWo+i+8419b1jgxUcp8W
pTUoLMUbQeHCsoA7CpKa1B8IoxpmYDPIyIgpvac725kEEJza4Zwk9lt6kCR/OE+2t6XOU2nxtKlK
6J5y1m0jwTl/a3LXda4p1oj3xch2SR557mab4vOVQ6qgKetzt+7E8JVe/uG2nUCipoymydKaR8ic
IESBlF1xtfuxvMSIb90uPhqnSNWJAANyHFsEZvo+znW1dEovvSBF6dfvrzPe49tjU8CK3LeF4WCJ
koP7FgHYyl0EdowRV75B3nq61pqfVH23ARp2Zd0jcx2vG8eXoyFgjCTybebzx/Cjg5G7Crioa2Ks
+3DIbnnA0QGacj64Sz8X5Q4Baqq6H3o0WDML4Sm3n9jjeVBDg/6UcF+62hqx2ZYTFzoiydDU64PX
xmAyknMjymm2JbIhVzo3XFR8/73s7nCU1EfmIB0yKOgd6kD+q3n13qYiqGQWQ3rbDJypLxqEsIuw
be01KACpexotaNb3p6AN4EvOzg/UglZJzlSHT4HiRs/nVDQ1ptbso/g9fQEm6MR+/rZdXsHKUKvC
GDL257Cmg3DknN3fJHpKf0F5LFxPG5tU7jl9I0DRB62ELuxMG7fxhZx8Ohcujq4VmCSlgLea8t+5
dIpkVzJjMrn6RFyhUZ156x51GctDEfvi2exJybmrk7YAB04BZHrGtSpamQwEIMwX90TtHPY11LsN
m2v08g1Fuda5jMrR1C6JcA5tYlRC/FoPlHMyc/8Ro30Gk1CwFo85nmTKkLRqtvuO3DjOjMGE8AeH
P0+S7eca4uuETw+PuYSpTFnmJ3Bnf6BGciUBBc4zP+StEhYpYSEyHzReYoHp4oRV5IUGVawQZ5VK
IV4EK2qIg8EesvhUSN1EqBrqofi6c8/nNI67raYYMmUddGfzu30vcjXPuektJ9I3WYJGCmQbbe5f
wL7ukxyylKzFRSJbIjCKEwfxJv5VSHrYGiV+es4JI8WG3bYSfPk735NFt2bE8uiRD33XF30l1imP
ORaZCnh7SadWJ8hSuOcok7PVBHgB6elDhXidQ5AmHpUo+a7iDwCV5/IbVTn306ErtYjDQAP9YB5K
I/oFdv9ylTw9DzFt3ARaNVmvXXMQ0G9AskHogtjwr/UweoUolhLDXxlAd83t9AqRcv85PZP9D3Bk
xMDTC5iGksguwx4935onoN8/GkIAHWirs7ghhBcwUxIncs7GCjg0DcbB8iWXx6O4kgZ/PYGAunJL
2DuycztwlQHfrIidn89S8OIcuILHfRHzks0OC4sA4UtfiLpa4BrdypB3YFRK1+BNR0ghN395b5Ni
JcxUs7TRuTQMW+HLSb29nxJ5EAhKqU36Gy8JJxXuH8b0Gqc9Aqi8jq+dRnAnOK1QOKg/IJTsGDiR
tkaAAvyCtUS2f3G5dv2rDr85S9jknCfQm8e7cSZpim/SJeYkXPbJj9gO80b/hFi5COO6I2aqJ6OI
vt1lYpLQBZ+Ur2o0/QScSutCM1cTGRUncbiKDNlq8JlYZ8zMKLRNwDXvjtn84tozYJY9tMZvK07r
HuwwTColFlB4cpdIa3BNfKmLxmLX5fqMq3ov1XLlhK1IK/Al0A/VZyTEGI0hpoAl9eaiDkTGvhrR
hqKQA2dHdXqlxLzwbJ85mu0TIP67puQwqBfxJ6d7g/b8NSuaid3dgRnZL9mz6ahpAyGLN3jdhut7
w33bEWATHXrmACnrzVs72bDqZnM/J2MLDXc83bRt0aMOmxFIhvKLDyyD+iGxHevP+SDBQ4McZqAf
Ljj6AQhZ6G9nGXW8Js1wRB50DGa2Ndj6AcR0IS7yzWVqGsb2tsvaq/ySZC22oP4R7RY+SCbp7HIN
CAkPWHNfLTSE2lghkN3M6gSIzSuM00oq8XvVfkLySoBg7/F/s+Vhnq7unG+ua2WseWUe5toiX11L
ZcBd7lx5KE+3HIw/NxDdsx1awamkCfjFjhyd45tpyXZAC+Uhv2lJ0zSgoaou0sEZTiqht8nkajRj
WpYp2OvCXKT4m1AU6usi5D/iHlbkFQ+n6eiMs0agzKCj0zG67Q0XyKfe43eBuMZv8BFWBx+KQogB
hLSADbl9Up+w65l8zDXV0IZ2if9apcF/Rb+BorQwROwmAJ0yyP/2tUWiTSWZTwnTaI/qdXimwNaS
oiQNUCVQ4shu8yd3q42fxH6Gk/AsD2b5pfkE33ItcFCvaM0cZpFXN8POWKX0eYWT6dPLekiRjbu3
VQ70lwUpPhiYYHs0ORNiQlxe7BiM5QLoy0KANuU1zGstfDMZJsHXQEW+AaokTSqzferTfuEylo+K
D5WFdpoZfpLR7PlDa6FxjUFYPcEMkyCOfFfb3GD7TekVPqUbelq4soo82aqb0YWAFmJTltXFDQmy
B61fy8Nnsy3oFYdp5Sfu0UP3GHGllVW6QWN4bKNlw1ENnWgowGTyZVV2hsR4+qBd8ym2lZF6Pk6J
iVWzm2uETfoJP62V+yDmzi4SzAc+ycM/VQj9YgxiKQkPczkPXHa0vjczAMzyrHbC7EuLPp891vb+
PHxHRT2lFiNYHp5vF7gUnDbrBXuA7I+64hFkpNNDxeW277tClEZG8kQ/2Y0dd7jyrahopxJP5Rnu
70lyL/1kh92guNaphWPoI6f5p4rM0Dnb7c7DdV4+E3++N0FV+YAVhr2SCEtr6wLcR8VO5Xctg30H
LylVzQtD8atlti+KPj9LlYnIU4gLetHZHgNh83yRRl4+ytjA6XFFeoHS9MED7jh+kDAHzWat3Q0X
V7xqCGeqp3uj0oMKVU677387CIww9nGHGUzK5CV0cIvCH97XzecifpL7jaA/KbBpDFsFSckE7jgH
UTt7UhfD1MmoLxwaBx7Ur3AKsQsk2Gm6VWv27ygj5tC2NYMKz3cDKeAGfbxvh+VRUtcla8AVNXt6
pkDvmUtjVOZKFwp/7ygnOx/o8Ll3Y/fXSMSUTbC0XbWUuF+ZX1rdumltcyJxDE4kQFOK795mfRQU
cGNVTmxrQR9ElT21PpTQtO4NGJtgeJlnf6T0tMvQzJMqy0MBCvhwLg4wUa4oQ/AsT1AvETF86NZq
5qzkZakxxHynBFslhvzR4r04IOSpEOQrPR5Fd3kSDjO97BQqUu3lNiEJBzKXKPzQh+3GyHFxC0AH
/7W0FKYNrdljRLF+VklmWHFdVvNIqqWArap8sPHx39atHMM366p6ehjNWwlXyV0nSR29tZ9vt7We
N9/hTbiLgLOPqA2hQZqFIxBMd4HQLG+jUs9qfLgM6+rRJBJLkrzvDpqI2y7F+vJ/Ho9aXuQYdfQ7
lJqSNQM6I6tvUwDeHZnMMEUYxkQEwqoaminrZ2VYaT34qt2vVN6s5n+ZXDpOjQ8X2y5XpyuK23rK
Mtt3lFlERi5m5lFWezcjYKH6L67b35MlLjOf9PJ8VtWmjmwMI3o0zjqcEcZP/Bms16xiFo6Tmdla
6h5i96ztUvwPipYdSOtAU74mZNFhGGzP5Fitrs+zIjoSHlPCe0wcNVZqIGL99BXi7pvbAtKIMJ5p
iV8dJCK2b1N8G6PtXJHDLVtPKzIhhlS9ddAC5vMsTtHxlrvBT6IoK+9lgHrCi4HHYel2mTeMj2vQ
dwm/ENnxpiQmCDcrhDnB4T6bnKFFmRxncAiCPXEKi4EnCACAjnZ18Y7BcR3vb09uJ1KxNQ9lZPN3
n0qftQ+nBkALbDU5XpbzRDsei8wMh08zLEq34JnzPXPZZphmEt7tjtTTCIcpbBhSHR+j/oH2roWU
4miydG0oHvpXWlQD36gnyXgzDkxHXV/YpUAKDz6CQ33uk+RlTxK3xXZ6UpaFSPkx8n6lGzPOUw0O
nxjWcba7Cs2PEoTrs0bNxQmkiKwTN7buFhxZULzgT6hMhuSv8QR2YQ/U+ba6gp6ocBJ8UeWaIUMz
dtzUjonPgYFp+JCp6M2yqKJ7XQLi7wxUdGRj7SLMd94ipGUYFau9YDc8KWRMnsVDH+IXnQ17lDzO
cX7e1KfKti0dg+OIUlz7Gf1G9pOyAegRZaBvWIvtLIoy8sSyY1FaJpiNH6GG4OgxtPcn/38N2pfi
WaqXWYWHKY9pZRLyt9rEKxpXXMzy9LuhNXjrF4lrieyQuFJT0+hH0AiSod0eYMC2V5wMCoT42hXb
LD8vOZkSdjQGtLYBfgJwXbJ3knMEKEtwHf94Yaj63Wn63Fr8cBaTqXO8eUH/u6oRA+wNH5L84kNC
zs9JP6i/1jGEouoPkFBn4zM3vn1s6ty0kkLMW1x9hrhTx6PVrorfqMcF1x6gB3XDj71kIDCQ/U4x
17KxPSn17vZ4LMbkm9C0lMRrgHA5MI8ecjp+C3BiIrGr8GKefhxEJQB6Do85H/7ZZxdUib5ltDWt
r0/Oo6YbSa09adbhwwNNbOzjjAHVOqxv/AnyGLWY+Pf4UUykR8LWoqKECNUQ9S9Wg7gPHhHHaFHk
gXzMScs5l+9IhJRfD6VU3V99L+BviAYWHouaA/jC7PhNz7qKZAOO5WPS3WA9AZh3lOxdFmiBxY4T
IM+0ASmvmroer8aEvrqhwlTY7Z+iDKw7Jh6hemdCDjgiBiWGEQebfLWj8mNw/vjWupmXidFF2gjj
a2nFJy7Tyvj82U2dH8xQdu/8wdUki1AbEv0mr9xTxoObZSY6VPSoUNGGPScDxwOQ0MNWcIEUvHyt
GdvoBWJxOW3CAmVtbW0fazXjenU39Z78w7ytzG+dvgKvkm1wVBSAYbWQKDuGhiYwRZ0BmQBAGm57
6hS6ThoTZYw4jRpn/ZtOSoQtskM0Nwa1o2yAwKNhGij2SgY67psf7k6NbtF0tUS5aIsombQmRz/z
OyaM8tsNHhZC2dXm/0e12zgrJECsmryBE76pjmdis1/YIKHAtWJ5q2hsTuD+u/bHM9NPYwfwuGKz
KjU8Ef0nKZdzN2n3H2RjAph9sUTv9eXSApl4zDLRdm1lfK5NU3dYQ1EioUkVVNfACsLdqjYkcbe3
vSo+nrbQKPtc1X8JpfNhDeGzPtVCBGqofMC4Bj/SyKMUMsBJE4wRBo99yGo8YwY1hxJRni/ADwjX
RniF1Ly7EB8cmAQ5jCYkGCQfAZkvKlF9+B/e3JsRT6hhl+SyHowxHAlFDtsYwHYU+aSzx1FGZNyK
a441BVZQuoxSKyu7WyMdvFSYD+WirPrXd0+4OxqHBoYC8lDJQz+9Ntp2ykyaKMzzap4Ivg606CSu
wOhHJwJPecDfaPDE9skhfQcut+k9yqkES2otafJb0Y8ybFRn/q+GiEb58ld6Ss8w/V9QSAv0r1Ec
Lkm9kpqghdIBJHIE8vIHxSdS8wlATynIwZWJtC0fNgksr53wqsnH++JumxN8qnGBH+VgwqHDmN/c
Z7lYV9olx0fWmVesIJqZLB9JbzR3LmZQd4rshqcDN0f2G7RRnaZBLIIzB2ipbrt7+pgY0+KrEgac
uJaY93s+Posu+aNvjjVcdUS5xbR2wyfBzUS7AFXE7wDXTmgi9kdqyEVMNevgoty8VZ/E6CJKEpxm
Y29GjEjTLa0rZyXPavHbxyNLNQ4x/5GgbvE+PgcmAu1XACCgZKg99tNmhRtg0nhO8oooq+WvW19m
TMotKcrxMTjjPn7Lj/ct2mkp/WfYzN4YYA12HiJzo5Va5p00bF4KK+HQFJsue0fL0bx8SCs38GhK
McDRNfwkINuSr58BfnNk4B7Wxl4YlQfVBtFq7Mgzelors3YRYDvTY/a1Ip+qekYo+ksYEkaZlKAx
1nkkjdwlRYRsB/qW3+Ezs7uIno/WVUjCtZGv3YFfJBymTriaZMx68e4jJj1llk87jS3QgxewD9IN
pI3ZGCVZMahi+b/UbGvuzhuJD+vC9xSpekApnE2lueFjyldIGMRSjI3ugED0smqK4VmPnfiYt63J
q+BFeDy0aCYcnbRtXupwGwXXfaB+h5851HBuItpp632BKfpWg+QYmvcNlZpR2mPr/o6lFe4f8KrL
bMJhwfKH2L9/Kr/527TAW7Y/UCbVknD6OGZU310o65NUBI4CeY5Qjky6L5JbpN2Ex6sVNfV3Nfjm
scGsdYidpi3BJqKHMSUYzTsha6jTbeGUL1512vqUfOAJ1l1ZxHr2JCekEPuvx0kjg1SG40Bd/XsX
IAln4S+F7oo9uruT9+aovx3XO2cueaGnutondG2TjGMs8lgo31GDuk0xLyW36WWAABgxay4gizNW
9/7Vzu8OHwFuxrapTLtRqFemnBpzw/3/SKqI2Fy8ttUBESGtfJvJ/e3juh+wrULudyUurX/FmhXU
+gGyoK0NXzQdUsTZGpnmxTETVASVjOf212HOYz458GW0xKYFnOnIoK5K/1IZFtWuwAGrc3QXIgd2
SL9TFAkGA73odvEc+oFSGapuYqYLfH1duRFo0nvVdpWtURBknXgFrrCWi09gA5DzNAuaH5HT8VRV
B7aaIgeDI36Sj7GwCNAC5crVAneClvvNH4b71XfExdxl98BEDR/JkklyNUwsA9EldBF58Wc536AD
mlJ5vztvDaJiQjD9/fhWJPLEWHl0+pDsJeIIKkaXkybrpUk0hcaGxLh8WHtto0JUNhnu9H1LEb8U
i1aFJeeth+CTk0o7c/e5YtTt9giQQf/MEouPq0kslohNFZItFZIOdUPyFnqyu2iOi3dHZL8Ejhdv
KAwKfozM25xPyBrXCsRp8FFrGcoGNIJ4O1oK0Trt3Tmf0+8cOGyKCdxPXyULWiv2sygJm2Yw30ak
XpKmjfbDXivGLDi2z0HodMxYVjef/peJqGm2wpbPIABpYi5a/Yul1cFqdU7Z12pi/czRV1Vu+Ruq
uvx4JIZejb7c2XuEmjb21qbBKWXiINlsjtnWKPSuRmBeTdWIhic9LokrcCi1nHdra0y8iZlbI9eD
zcM5oZKIZFfSZyo4LAczUaNAYT/pJPkEa0rTdxSjPYBw/eUUs1VgnFqf9WF7DlaIIeHKHLqRqyMa
A1L+ReTPUqFmFhwabq8808ZNVFilrnZJBtGqADZmxSG8oIfe2/9abO0orZ37OSC+vmP33jNNgmER
T4/2z1UNpTEXf73Tlh9U+rYsokywHx0zldw362WaEEq2MOBQYf3MxXK/Yx7QJT48yQXzR0r4nY1a
FPDcyC2so4IyWUuXOcxDxki7wg/iKe7tCikxtXmpag6toZej7/SiRLUwaqaiI4skZb+GEPLOc6it
lzZyZeYJ04ud3zFQSKuyDfhkGOrAo60baw39j5vID4US8wdDGCqrJdRQ5p7+2CT/rzwiNY1ln+1/
JUvS6FG33IAbG3iZPyhYKyiaD+yXWuQk9jx0x8w5qNavF4FIGK0rq7ZjD3QMG+YQ1eTyNUWdKQ9+
nmFqwQQgHTZjR3ejxyFS4B9T7rExf79q1s4kP00Tl85waT6uUaazc8uJY/lmvEryUlZszWbHwJja
xCad//TKBgSD0Ahd0rAWqqNwT/jXD+IVNJI+rsfD28BtLgPmxBj7BjJhtm3uuAhRrRzB/2VNDIRz
4Ri1d5mV5vcKgpYE+qnaCui2QuD0CinPMNWPoqGpGNWTzhpioi+DLL1fS/HmeSNuc4zYl/oTGwgE
d7S+YwsCinmz/ilwO8UhElgadaW77XZpnCxMb9Inul54MIvrgulggYBYN/BPD6Qyyfh4AVly3veY
6Il+zu7VD3ZLA3junQPwuXj39LSasB3b/19tkUo2HAhMc5JeLEehzMsdCCJwL95bav35HgwEz/vt
PKqe5u/a+aUICNfax+9ZL6KczkobaDZBbPa/zGuelz/dZD5q74vosSD5JIvMAD03Xym2VwPCab70
wQFTyDPVZssKJbLq2yNu/rRigoculcGgaJiAi/Zjn55ReUyMkYaoU5Ss57lO2PuypVs0RnLwFI5L
ydrpimA7AetJpS+sYMJBHkPuVtypchvkjU07ImybWnL4GrUAyoVGY5ejp4yvZtcSES7aRIM0KGll
QR0PcZN7+NxRefdj669oFQrh4zoIoiasqd2RBS0iGEHZQ0Xai9VTsVZ1jvewGG9ZaNfhLxY77S/V
xZGMCCnvBN9oCmOFczoV/l5MUyo8CintmCbO1QtLx7sH72nMzUXNaj/OYd0qJoJDwWCveBlbfk2m
cb4Y7x1zH+9cMYTebDS1p1FJsol9h4GPUWWK0Yhzcc2JViI1yg7o7HdUuFjJ70wAhDO51hz6Z+WE
RUagPrNqsfOju319M1sIbvjIeyKC1WNYHHTTNMenad133pvXzbHuSznj+7JH86R9Mw+QKiQotrlv
QtdzzqFw3ch0IEVkcWQUxSLBm0vN3RNZfAW+7uLXeGv6LqyfaodVTdTJM7e0muDo3L29nLlqzkhU
A9KSEf6uEcusHbV/V4MRxJgDt+Vgz+FaW+fw1NRHAbZyw4rrEyfrRr3rvK0LnfuT9rYwnZIJfpkb
zQ0/yrLuSwlh0xTPeNlBapWU0Zot3lJ3/9xNqrnYMoQ3vXi5iarYmi7yOaBHApfp8OEwvbexZT5Y
NCdLs95UV8firijVWJ9JoNahNODLwDIDVwXKgCV1Aa8lYogGAmCvUgkhKBlaxGESqtW8+JDVyUJc
F4zE1Mwluh2GDMpGOS2hrKR5oHZxcHFboFUOq4zFQ/Ub62TA1OkeJA/YAfrKckUoI0rT4YqL77O0
+WwKO3YqR+fGkbq1oVp1ZPVJSu8UZKdm+Yc4mDJyUZvJPqy1azgAtMVfQSCzBtxrVtZfiN9dZtF7
pjstDp1Hvjos3QlWA7pmaeWZT1i+fVseICToYjtashQT6nid8IztxPqVfvH7GTb3iNt5naC5pFgw
z3pMYBRA+DYTGbSQLLCKlt1QeCYFXB0Wops5UlLlB0VthzIiXSCSgZw4cmWQbiaV+14Ju6b8azv/
ymgBsuaELvg5LgrhM+BIyBlF9NhES8gwme9g1DzuENtxlLveff9mvpzhdHTlTxrO2mQvvMU2cgPj
kCZBVcixCaTmmQIMV6N+XwLoZx/zg1sxgim6ar/10nhkn00JgHe/TYvaqtA+HiWB7OpEb8j/fExD
sqHC/CuphHLOdQGt8UL1ePFyLzIVeP8y8iUi4e5AoKx2NW+6QJKCK/N/t+sT8u1aNfAWptdbIme0
DCdAG6YIPInKMfQCwlesEKJfTSvjQoI1XytbG3f7fcAAZh4cvg5MqMMiCOkN20NWxIbcrY/SfDm4
xjPBQQVGtjD3hO5SUEw5PJZ7q/+foFesWynGkVbIsMR+NvSbcLOWEJCKe0v393jXIXybsJommUXt
5BHLNBUrkijlkTs0A306p9ZKD4CRUuXTIRDZQ5kXVCTWJ7oaRfRjKcjKlCQd0gxMsmubdY2OAZm5
Cn3cwmdveZm540Gcxif+wBJduS/wU+a9qS8va1MhSFlz31UzITdFWBS4lHVQNjq8YYUmEX92Z4dF
59E+FRRxneRxBMco4Ix8icBREtm5h/d6c/FJIAHoXNTg7FUmEsvqAb/ulO9v/1DVZuCoNmQc9wAK
NikeewhuPWe8CeSyxgODp4Iy/IzvJaVlJR6yJht1wMeTeiP8EWAPlmXbg6anKTOKR9iilTMmBA9l
WpufQj4xxhxtXW0ZAGjdD/UvmidMppPjGmsG03HMVseUYgb4Nyk5vqePOvAXK2ol097uEL3LnUQt
G1g/D+/NFlFWmCP0/dJeIfpDc7OnmCU2V0wYxytJMduqqGGmFD3VZoNy+fJacuR7Ty1bJIPwtTpK
fxa899Jseh4yFqJCsTa2qxBUucEsuutyTd4hH8peKoZanNhcv3Vs1GEd5ANO7bFrTjEFb7cvE9K0
GH2FmkCDPTHDhaxiHI0bcmohlUPte41q7cOhBJfkfkcis3A6y6JqilYjGAoQLixnI3aGM0Y9QFdt
gtrq4wkJwFY5DGHR50mosWfupmwwuDOgwSS90lY8CcxaOH2H89L+kfaPxAu697OVve6P7tiUswWR
qfZ3+UV6dSz27Vj7d4qLdsdDh1Mp0zqWFxuDmfoN8lwFO6CoSI6fTA25FWF5LPAu+22ZzqVWPwc6
mLKBBvKmeWZydVVo+rFAmBa8GfHELY4BlJ69kx4C18nciForWWHo9Z/ADqcYN32eRqQDIgnXzDZO
pFvTYe7lEeO7YFW0JC6y2pK4YhtmnWwlhuWqoNq2LUeDf/ECNp0Z3zz1MQDzecjpc6g7UueyQ9yP
4bogDUt/FRxEIpyoy50P+p3NKl8XK5FeI7xRBt9OzQYrV9j9zzb1UnMMsfzU4iLF2UeWSYXOiHf+
j75m1zmVsu6ByVtbN+RYfCQFUr3bgpiP/Kk1Ni3aoV6YouSdNJnC05QDb2W81MAzOGDX+Xs5xxIp
pVxdKtiXegK7R0qBUBKHA8CBhv1ICzR5LSRd1+ptuT6sSq3WwwC/MVGppKc/pmD+WQ2tjzMmJ9Xi
fGpBeWyPyVmcDEXFMTN0VnD0hAUacuZdNM82GzXKIV0nPuiO5MFZ0AS6vzrGobg3tOUMhdF43h6A
cm9hYTJywFTm2cbIUKLepYZVYLROpTZ+qYZQqFmauYgAYyJPTRK0aiYEXKL3+eDEYPvr+wnJnXoL
c5z3PwcugOKZD8k7+FnvICCuJlBk45MuqrP1bDZw2Je3K//z30XSGju3aGppyNivWQuaJjDFsNd6
XOdgET/ynbfcP5K8uQ9GdyemhiTCKWKe/Rd64TGUDsKJhHhGylKnixZJDB/dmgZe3wfasKIPmLuv
SopJFlwqeup6g3bWiUzq0sSRGndYavlGu3Jn+iazDJjMqpRZ2VzX2Ad4FVT4bUZguUDe6lLvUiE3
jcQFQkd4NByXSpoZCuSXnlkWu+dtUzO+rhomscEz4tApwnfcl0f4MCdu17mMLWEvOIOYwnzsxfb6
cgYTovx6q34qRPAo11SgOm2WQv13PoA2fkrQMbHphZe0b4pJ2pOVQy4N2L0ZvgJAxReTiIcc9Gh5
MLF1Q0Svq03iEIiXC1k2kYOAnFxNFwfVrcrqh8tV2UPRcEX1BC6T4/qLlFbCueflElxcJr5bGxDH
EsqK7RcOmXWkUD7CfUT/6wzvS7GYdL0qIRYXS+lgZyKzouY2R+jSt1/bxO5qxDhwIa35cGskFYcB
mYV2gOY0BZApSsSMWSCL6zyeukXDxplySMFjB3p/ecIe8dGGRDag4X2qvWDpMPX0u2MxnD2tq7pq
0H2lyd69JuHpDirZQY3BS1vmeP00stYLeTfbufiXoYiWOZAeYQBwDDLrm/Ew6v5zSZt7Bd9kujll
5cltSwHWv7BSLKNHi/BwhEC4qFPXIH9ZhVx0FRTOksWQybpxt//548PX4Bvyspcli5wBUGTDtvB5
FmQxOc/4oMqLHyS3y084Ux98jzuVmJ9DejCFvjDxSsAqQrW4NojDMq5gLQQvNkdUlUpll2V1XBD+
GIbXDi96yXp3ccHYxYpYrhQb3/VqdP8blpb2fmxSIb2/TQvgTliK5tG4gP4QohmmTwzlZtQeQSFR
QFVM1UFW9txiZOBn2645zo7clJIn46kh30533A0NUjX6X7xRLUPCTartjSLG+k2sLIHPUApCB6xs
rG48/o7KYSXsTnQ6fjn+ijt5x9uIk/Sek5BeOE9HVqS8ctHrjQJsAhOST6onBfESnaSSixw3fy1p
BadmFWfptHRwA5fuau/vlDavgDr32GEpZA6Oa2QPeLQsF/U54cF1xda2TNSDzJDpTqdHLJoCETi0
31o+Og6lY3CvlDVmHSfRjSJxs+NaQkhZnz2Zblva8/mqzcZvVyoJTBJQoDQHfIJ5TppXPBSi9Ou0
/W5Mlj+EvsTd1XhNXkN0BesvIUdWOnc+9CcoaC9ei84c3pAEX3V3uGLwwY6huUCyUmBo81dNd1RP
CnR6J8jXA8zrldU5WG5Rp+nSMA+vs4P7qQs+05tlKuz5kjZmxyH/UGGmk6SBj3bgAq3TK2PVkfZi
1shkDxR+cQPUT2XSShvw5mUan49Ow9wMrCI2TM46zIKrEhJ975IEQ8TGqokBZyC8RBqcZ4iHFVp1
uYp28DFAbnvTjOFP4MGyJbsobrwx+BttEY9Dy67UHrCXPolGgTcrhVTrODhl3Js+kYNeIVy/ZKVA
RxYBB8o09s4qx0/y23yWCv/i82pc2I1+2IkH0fAwRrqPhqvNSDhIeED0M7AOUN/5gu26Rq0qrkN7
Dgdx8xDcM2tvPl/CE4faiCfFXHqY1De2cp2yekLXXIKvygzBdCPdad0NJ7LRg0p9Ye6dfGnhuapK
BwLg3CJp+ppFDLNpZt4N9DSDuUTxz/Wmt8gZT1ve8CXEsQUBYAGA9LRcKusX4M3GJDHqH+U8sF3d
d+oeNOwPjkq83uFy7bB7c+VXFKQdAtmf67TrP1OmHLGaZwWNzwbDJyi1uPCPJeGkKF3nyUptL0YN
3REFBdLzB144qhlcv9zXqaVnJkMsCNneZnWdxppPWgxGlcARtVTGBG1c9ibLKTKFMpozQT603F6G
qY6uaDKV1j8vB3wcMIh+ulfKKqrlbBdxdmWyhT8pL04FLsQC8Or/VlX/0Y1CfgWh64D2RBEDD+/g
D4XYNqEnmBlSyrQNGIjYFgO+xZdXIRlRmMlJ40BGFnmM9H4BBK2MpQFS0V8zN0yCLl8sP8P9zz6G
LH6x29B6CegzlFMrh6rJjL2dIm1zSarxun83f/83RUNo3rfz+sKH0hF3vTQglD3QZWl383ned401
uJ3h38U4MBp3nuW1uyMnRLUlw7WSp6sJp6kfn+LTW3RLglMqriN1EvO8MZVDGBWXg0FmsJ2wa944
S8DxAyuSMXrmCrsaXECjLW1FJl/eP3Wrnj9A81onDm+xLfJj3N0TKqCLqE8p4WaSaHh43nuYeqZb
zj9A2U6FbBDSQ8SMVhz2QcIyBNwDkvyIcgLGnRX2wHT5y1SvuaqF8hyo6KRSTsAcOHwSPhfnhcFo
mX9sX/kVhuGdSj/KNYtEHIq37zI4OuXj87gjKG+j4EOdOrm02RbWBJKZIvYQx7Lf5aKyWxdwGS9C
MbP0jRdqt7G7iUFGD4Iiube6P3IpfO4oood28AEvQ8tD0JX+zX+R05VA+vZgUGltQ4mAhCechkc2
RrISBq3ovkiTu5EBlcjYf5a412eOQp2QxT4Pw0nUbzKCQKpDoNFqbl2phrA4/0YOPz6URmLyJNdj
bhrB+sb/9OFJOCzHcFixkm6y2QAAFby03DLLzqUftzp4Cuml0ot8SM/rqwusF1X+wRCo3odnkD5O
0861+BlwyAbmlJ5G9dzkbKiRkz8e6l0nQTP44R4x0viZ/wXHJHwsI1GjdoMt11WHZQnKkQaCQlta
YA6LQQ14fZuF6tXbU4u6dgqsjlaSbe9Jn2Ybcg2xQolValaxrb5qZnbQSCyAgHwCKZwJsK9wHKG7
ryfSRIvUCZDo+iqozmPBdFhtZNqQZ3TU/N2LikbICi3e68oSRjDWJu/aKYc049hatgVn/vsChp/h
bnr7DIg/YHfsAuPA4OeLgtyiaCksGWsMaed4odLog7GBxoPRuj0MH3R5jGadjdDPOvrqD9s9ftjb
LG/bsE5E9DmGxk1Kdzhu1gAMsD0Vb4NIHNJC5r8dMaw59ZqZlG8CQF00pP2dxtiuroonOCqy7jtB
Ulc8vjFAMEILgxtJjKzp/9O86jdBGF5aosfVxd7AKlersBrz476wZu1u9BFu6YxzmKjovNPaNUUd
C4PZ3JAiCDdwr57NJua2pRiMpjcLyufqh9zymMK87tC8qHSH/yO4LMWVlCoSNgK9Z+8ll/1t0fGU
ihk9yUYBgJu0n4N5Jy6/f1nhwlslG4jPnycPbqLbmqrqn7SatEZV1RlApVuOX+zX3qUcO8ZcatS1
4GAbml5g21jwg3hu19zi9SXo58eIU+fx4tageYpeK4kxrp43cnGerw7VDp4AI0LtPtSqxcHGTmEq
yAE3vwKt6wZgnAmkBFuMDRo76xr2Wh8uEePgKBNCegE+PZldlCV4tXWaRj0ZWTMCcfbhUHTSwqDl
QS7O/O5/3tqZHkEFbJnDuSjyEkSzn/Y6gNl5YB9zJEpD02f0Js/ae2NCJ7+wWmsT2BfGOmdn8KGz
p7/o71qPcWRE5YXLYenqp38kFo9CSKFeA/Ko9LfKTKsq/VTUCjAtVBSoPUjpzoxYjjP8r6FBnNup
1q4H4xgo55naIoL8FTaQrg2wHaw+STwPsCsM3p1y080rKIK+iqT94fGKyTJDbz6jvs/4nOBFVHW9
XkdiqlN3qsBOc6cH4L4r/Vr1HdthNrTGbOuVplJSQ0vMucJCKdAbgNljmEj8iwGw/LdGlOGc63hd
bHX+823AcgrIe7whRE0LG2s9dPavtkGj5wG+L3jqg4TnW90SFE0SYYCYX9t5AQds3TR9NuzoR2RY
H9rZPXLDM+LbdfxNIUq2M1pNUM3A9+3Q9eMRydrU8ci5kBBHUEdugTFj/zo0wZZHO5VEOF8ubCIk
5nJLuv7yQpW6l8Hnn2WomCwM+WPMGDUGCETlsDdZSAOXLocY7CxsML/fnVhJf9hD0z+1nWBYdoRh
4Ge0TKTzB3dSQUVVxzWMMTBMOkRiWFgDOZGXVmEVpGo1IcYKf8hmvWDJWiHG6cEW38Z66rvPrTo5
4qGXkAet8liv7otR+0LZS2N1IG/07+1osEZj4b8I30g09w9xd8/Yg9yj9iATIfo7Tt15Y0oi5fWX
jf3obqoDprcUe4Lw/R+n6992RTZ4fFmStgWMQzd+rfBllmv76gZ9rbYUCtjirAi37HkRP91NHwNx
VSaFsMwuOSiBRj51KjBVG8DCB03Sg77sNd6D8rz1hKMy6iAd6v+ZlhlwyGsi2YGjwFYb8QEMfVSu
0fYXftsMFq8wRmKZoI7RGTGaCQvqwS4WZzvu7MA7VVUFMhtFoIRwfKcFRQun7vD4sdhbvjURtBqu
DP+Nc2RNTn5WVGun8MkH/+4AEAslYKa6CIfO8Cez7uKNk4CiQlG5JnNqefZymbEuWN/MnVnH6IoZ
9X5e7p8ZvVCNW6EF26XBCV8yg5eVqA7d5GQVwZgJ8KRn+U2nB359DWM6/BNRVmEOP7/M1dL3oqBw
XBncBZ6WT0IDMNNztdLz1orye47FppMStx7v7BrGmRLHs4ZJStaFHRinWs2cAW+OqS7AhS7tr3Qd
XCB+KBm7JSkDqiXLmGmXQLgc2XM4cHMjyVZ0qBiOqEHplJkf/qUBsk/yMs5Uy/KTbo0oKZ5MkKQ4
VVCTyyN9ixFDeu3CIFYUVhV9/X4gTCE+rlKKH6rBeFYoJfpaSzNQP0WGOxnduc8/Z+z1hGGVUyie
z7T5MFCMDvsZps9LAYDJZD1rAVk+l694JfH/o9xpzVLv0gfUiRGnfL/+UO4UkIo57nLCZi8f0+yO
HYU0sClwFN60hrh3FGwWNcT/Ikp0J4en+3U5ZhAiwHFPzOS0MXM4+gObYjJiq6AN6+zjxGLg+nMJ
6oukBUwFDINfbc6onkZFPqDP+TeRZ4sOqvwS+bgmvJzjf83EePtaRhegSyLQxMKPllirONFoNhTX
pT2Sq5e2y+4WwB7sJaneRFd67US5sAG70J7YIOa4McZhFZOCe1gUm3JrPQ5vEPKf7/wkjRJi4Hvo
LZQ3irUkicOc0Km6C4VtBZ+00FVtW23sGsEHlAHYnDPn5VROaQnpTIoHOWs5aPrJm8zSGlH3bTcO
o7sNOLqRMInOFLyXGOs2xfngRahoIaoslU7HvD3Npb8VOtytyiWNiibD3X/gFoX4PBAXnmoXmPT0
ENBOQjuYo4lpOGR++LPcLR5ZeNSjySih9W770MpbS30auu/MSmfhJBF7LShoYm3RB1iHLxG+H904
C22tUsJ7ejiao2PVDKUXprnH1CWLSRoM3w5uPZaD/cl++/OW5hkioiPfqfApvg1/Vu2JRBCh03zc
KFqoEtzvFxNOhDe0ZldGWfYcyakgGRd7XZU3LfWwdYBd9s+SyHzZpD0nik6z0+y9FLGyB0vJ/fYc
fqfe7nZpq2Ke/WbJ71zXz+vBDhHen0K8uQ1hYyffc99XuJ5l4uoZAzAY+cVlcjIPHG88Oxym57ov
5c7SCxdSt3WrApZYFil+woVFSAVrcLQbcBJtg3zQndwkmf07jcDWcStNafbho8nKI5NSArPW6lyV
1F8HUYZWH3QVMYhLLJV/FGQ/X0+M39LqF5CMbKvihFYCluDS1zebVUdFVnEGrItXp94GYjwfMg1x
guonJLUik/FYaOF1F8D8xTqCA7NDcdOP9IjwENWX/CdO3f7HN3u0wlDKkAU2XnjoZvchWikjgYma
+kZVDbWM3Dm92tkdhyD3sHKIXtw03qvo4QRUi3Xy2+h4cpJj5P+RqzR7pGeE1WFApJHzb0k4yKaA
WQ0pUahZj6wae5ETv2uETmgoA8I5ddjRNCFGGo7H9RRgKDcnizihRruV1Qkre9WGtfnqXQ2HZs+F
D6Lh1q9xn0QWlLZjplec6VUsRktEUMAJ9WwT5KdUkY5AoZ0X1+ADI+kis6eZoF3YWuL3W7ewPf97
HN/0f+rMyTDZrtnmNhAeT2Ug8dtNiV90/LNdhu5JrsDHfrEOAJCjEctALdjUiwcifSXXCsW7GA1I
DqH/TfRzJgE543XsplRtCBXqJjqDtGjBC/T29P8VPH5TNs34w1ZD7eeIrmDSzEDiASOYViGwa4/6
tx24J+2Wn1ZOXRFn0G7fQM3/xo3wEejfx0MSyqSHFJrXPdfgktM4+8DLCZsgQbzCKoQEWv62Wl57
ulMPcdt5ge679+DBUT01iPeFwQk3fCwbLTaz49eDciGNKmX/BWpp2oXxmSX2yLrONnAAfHDEJcd9
G4YqI+X13L3/cH8APp3xhQkaJ1bbuEOFbT338xFBEHyuWBJxjQ01hUfadGUCrMjOQa2ApZTzWyjZ
IYOSJJ1Wm3KYYihFjjnUzwUubX7UMFPnZVOAJJ0yqthQg2evB0zFqYaCCRjeOCRhNc4vEgiA9AtA
WhFZ9oZPV9rYk7VDScWZ2s761TK0n+Axb0xWORYlsgWF6wn4vWjihobc1afa0FQPT5tfMBBAn+2m
69EgcFnTmRIjYinxaCMYUIEXFUWh4kM3c0FYyJjTIsh5vvMXXuCASCAL3H316JvMY2WN3m0vt0Ky
Y4GBL0e7qGjxde2jJ6jWL9OI3Ekr6lBrOnvJseslFohHW43W523ibNYPsU472TPzScP3KjORSXNF
m3YlQ3TYkVEqSjflU4oBk6c/5DWv24UGsdFByS4ojOymiV4L72Cf1jW0JZs6ucBfkdatZWt3ZPOj
HM7zWT9WPK3JRjrM5TGL2UTSg8bSRi+Yo7+Sb2lzvGY9Hfqhnrf+ccQ360L97ppDl+5yyGCj8GsV
yjUj88mF1QOFRjRCFKgU7V2EN8A6WIhBF69ulug3+R15rzzwmGIr+QHsFA7dXfQznGzM5f+W5nOf
ZXzmHdDy2Uan67amoDAX4sLJpKL0v5PlxOn9w68fjnhav235FBYKJ+OGLpcv6nKi8O/yA3ps53US
RaiXVdHgRl13457/yzQ6UfUIYL0lJm9YcRT286vsi2D0CWJ5aouD/5Yc7t1AUDEJT9jf1Yv4ULiQ
SbWeeIUFvC+vkG38vV1RzqhKY78/HTvpfhLZ5KUqWgftcXr4f0jhf2UH0ThLJ2yd5fCwnXFvCwP7
LGbgDdzuxtfrKofwbbnap+U1uEZ1XtlHejgSxrY7VxP4izoILS77lwUoW37bxuhLBq6p31jRc7rE
abe9Ysd1Wsy/KXA9GAmAluTLbWcGpLNjTdpKQVGY9VfSJbbjFRlzANhuLc6uDhkoI7+pa0ezbVNb
9Xmo9JyGZD5vLtY9xZu00qm1/2aVPoOvzd/ZohJUF1RD78qNV7ECfvBZ4b40tfU2kN/ek781Of9M
UWhaLSm0ueLlMHwH/OjSgofJPXH/6filAX5wF4Blx45dmLYlfwnllztNbI9FQOcbS8y+hjSQARc/
8Eier6H3oY656y9QcwCZfTBpGaEfZfiHEA/gmzkjUXZuadeP3GB/MFaf1SCcF3/yldhLDeq5/++m
IuHoaVZ1ZVeTI5Suhkst8tW2EcBjtX9qtNrLFVtAMdIaEpYc1L0kkHisTvtL+9ZMmiEiZO+LsPJV
+OF5UeMVIKG5LBkJTkl3i5j5Gpu8UN66VSk4v1+ULMDrNHv+Ug7PvlRQsvr7ZEMUFNgW4K9U+9WT
N+POitrZlCcni/uPl1OJwuGgRFRT1vBK2r+eOG1jxsUTUpJS9PRTCLob4iwAsOYtb4Ir/+TbEZr4
Ngi+y9HVbfve4CS+NI0gnKL/kPxw2tFdIsVdBMLmPgtXiLZMuxuq4y6pCAkasoiz2eJO9dqGzg0W
rtZeTP8FSJ8909ujwZGBDclvSnhzGetrQDjPOIDz7pJprqJ3ObMGRvgeOyPflUuyQBvF0ChDIqJH
Ta+zRTYznWnd+x6ORs4fG9Pt6yss5s3TOhRsfk1xrv+PT07BtevX/BFjFc3SiMhdg4qUQfK4rziq
8yebDpoN57dyRM+Xq5+RmBKeDcKmgQl+RQOhCLoSJG3XhIBMv4yJ1jcB5QJQXR2ng/gG49qePhqH
NGfYJ4uId0xHecweplgd6note+C4wCqKbLYwG5S4otUXruxm3d7/6YL1yUzMvxSKlx4dH9dzCQym
U+gx3z5FEymySeaDJlhRDe1h9p3Ae8aA+1jA7n1oMIl1XZmj/5RZS/7Yf7sNi2zaO/Nk+fBLx83H
ADJ5RmGEdhMUuPE/0IrFM0KPRQTE87tJ1BOzTnxllAuiNDIm9hQGVKN4ezxeOF2MTItsuk0lolup
ksVReTlvR0HMaW+I2dXqRmKsS4MbnUyTfcxtdNfzJssZDiYzJYVQx7zKweyG/nHWfI0RN0q3nE1f
yhBXK0WPOa3PplvT+UpCAlS/+gQyjlNVc3XCcICJqHLkCwUwQzdqpRPsYgyGtDeW6Gwf/NJc6M8S
F8k6qT+C/khK/U4H8Nba/EvBRywKZsJ5Wj5rH4waOvUlqNoyuBPNTTKHhYAkZlar1oQ0H9XXBI8Z
VMuswFdlCheC2NM4WoLGlhWyNJNnEMuR/ysW9Rmmv3+x+JetEq+YyQjcf3Q7TtuMwTyIhqxd/QSK
zAhKXQYVYso5r4plM+RmVLsyE6QvYHhPOAzONw/ipGIcOK/zBlNyJLZiO8l1jmRs88x2k6rXPTcj
UF3VwCvzAje5WoCugVajRBQUaw0YwaKV/sdTM0kPnmBBrUIlETOinqsy8/DsaAoUY509S8bNkkIR
skpkLDMFt0ZcQljWDoaLijrpHAn/pbGmNOKtSyCpnMftApHQBvVy140gCbcYy+gcKogsefjf1HhD
hqGtmqRSg1CfUz47TzL7zyZ5OVDVlCLQ89C9DVI7G+3aIwdz+zJ8R3gBvVY/cozs3ch+8HhrPnct
vWhJwCR35TtmBIC3GtfbB15toa/b4XgTzOcCtV+MDzFCqe9jdq8crrmAeTpW4CStYHxi5MAhJppn
U3T9l9WBE/eakJa+QPVWobaBa0Q2jNiLczDRPG036Q3/mXehKYxAPLZl0jK005Z2Gjylouib/7il
5ZPbqh3z5a6fo5fG7wOXuCDtH/ytbXuCC6exzfWGYLCf9j1Wms7JSUVGZKxOWlw1Nq4fz6fGr1u0
tuyaPtq75t1KpxTr5adWY/8Fgo1+3omskhnKf3lleqYxRI8hFvd923DUNxd+oz4KpoAT+PCSciyY
mITgCsZApJOWyjbxY30/CiUyXzGJWi8bcKhZ+qlBNC0Wm1XBjKwfmIdsDlwAwp7mk2v1q9USygdn
zWEJ1T1+Oyg6PAbyyacNoPg57CwIBT073EHqucratj96NnsquqgxpBLZ0exOh8EyYbAOMY4jDaFr
AexvcJ1HOnMzpJ3b3KIQLyYEFspRlkcwtRAyw6eXDFguYUMRTqZb2eV3y6udEavbz+uoP4XwJ6w1
INnsXz0z+HC0BNbwA8eIFEB10UIkMjmF275FQBDVxA2q91Ce6ZSaHlVKXsewg7g/pYnHtFpHNGUS
ETb4qx1gRBYFMyTirDh3K83RnVrgtcNN2xCs+YUJxiPtzbOk9Dag0TDAoPjYueZmx+94gTvf1ixG
0LgKIQz9ThOWKV3CqhY+t2wpaZxRmz2pjRATPMExsYNtGD97ViqE69zPLxLO0TGltey90YeECBsh
LWK1eZXakJW3wDgcnr+O5PtNHVdqvhvMpLvIfI5q0LYxhrPKZ3UDLoBhL/eJTUsrAwEOA/lEAgyG
wlmrW+gfiJE5NRxn2x6Tp6ZEJnYvQSF60xugn6ZX6vepm0VyLRUF5fa+rHv2A7vMRCcEMVgQtwws
vPC04whjAMRPDAyT+CZUMN91yiYk9f7EKI72SSpPjk++2rbPQCb64vo6SGjD2yhbOI9pjuaq0YNK
k0z8+9Qz6pJZizOygAWK4ciwepIDW/K39iVzMKit2P5tR+XMBC5ZN04rYwUDfW+lYkD+UquS9xSW
m1DyMs04akiiOd5omveuajQc+jJDz8GqL87N7P2hKRK4QI5VODJ4y5ZZVCNIugmcwTZIMb6UkfVO
CRvBcBkR3HuV3Wf4jNaoKkGfI+sTAw5igCPwUNochlsAaWJq56QSR/pQZIi94tW5KhX8JeQJ4IOm
hbNxxhoPPvB7TDPVaq5GwkdxawfH/sVngBHot7atg5NJiy0c5DjW96+7xAureg5XAIpDHUGHOBjU
aE3TuamYcOM4JxV1GP52aUduHHbOdufrCvRADOmfKTsYTOhk3ZwInjPlN73lz6ZL/Fm3q0WtH5d3
QdRlwgbigLhEDc3ZDgutcIyDPqDQHmuZIQZi0KLFrv8z6ajgdTeSCJpZRlJTocYUxIxKNWireSvL
cZpheL0ylGinGLUPSjQDLBd7cc0XWfPCbF8GhP07XtXb1sVAbUtdbSCvguiAEt4PmJ8Mg3IrjJNd
zgIZHCqIhG79atSs0seObP57GyQtOHnrYytbUkpXn7pCVi9CdW8957k5OEtxozoTlPtDJbXYle0Q
nlRTvYiHvfkdk9GNUEOFRCpNb3laOHy655aAuw/6fvMJWB9uK6OVEOXezcR6yIMq5gX/C7m6xz+x
UYVl2QlcB25cK8wyddrEr+G6hT/wrNmwtPB4I0PKaqGOcc/6ssqnmRhRJ38/F9m0mTPe4y1bvrOi
b3l3iEKNLGSUy8sB+KwjwAbofKkWKDRk09RP1Psz15F+XDa3CJRqUa1yE1WbzJJAPfOPcHE1j5qU
cwiigPBFiKcBqmoNQkqdxVjMzJMpF/ct410yKMwoLUlNVzkiC06Pg/wgQL1cMPDaeUVHRzKXnI8s
+GLlcRET+3rvP1D6iVccF+aTP9pw/wN+vM5lOU4yzF2QLD2sFpSBVA/SuInkAZgIsVu5b05W9PFL
WmCQYS3H1K9IQBqObTDEd5hxos8ESB060kZEeBgwv1+4wwFAOdN97FmdwMd+Fk5zz8U7U7qf899C
CrWrLn/XANwDufP2d6UHtY3cWlcu+fmizozpG6rG4Z3gVmbnNFKizV3T4o4X/lTHtzdVESFJ+Lyh
joHm+u61i69EIuXPlPuCpAY6s6pHnRqLQIHgghSXPHDG66QQWu3s0UKcfeTWsDwA0naYqth0VWoQ
GUfs7kpCBEtMPvlNIGqgQmOjgO4NTsecdBY43UxbT21bwyZV5diWt7QMgVHuWfBlydnYm5I1OtRX
o3g0hDlMvnNJeBakWe7tc1NvUCjvXAfREcOM1v7cCg5wgrQLyOmN21jurxaZYsWsgR6hdPb7XTMj
Fn6kaPED0jRIoDJYnLQO0bUhFB9KzTjqz5Io58ZDmCoKYBBkQvDzelL3TxNIZqzk8kaV9ToiVoFJ
uKycN48ZAvRxveKMp3sVphkveS524XbwV4HLK8PngeoXAjc85WCw2ztoKm1ah8fmqCbJxp4GKOn7
Mmh2fe4mpOj4wO5gNBWZUV5OZmALXzLMl73BGmhjpJyz7735JVyJ1hcb6MhFBC4cfBiZ9XB3mx7e
r2/ZtRHHD3VD0xv5ZchO4mh9fMLiFvNBTWfP6wj8FN5H16oDU/JDQDq0JnXDmyi1x/M4104/Xi6e
JDYd/lgmCy/6KZZ+IUVYRzdxZkLQxPxvMVeOl7NJcQWW+FgICclV3jG/32rtn87gDYkxlnR7z25g
c9ztYDrs+nUI4bUZ2L91y5L3wk69IYXaEeNhIdre094CEaokP1kp3uKqlRsUHbnB+LUlFyE6GoxN
UW8ph9ELSPM92M2ET7k/nrX6PEgez9QhUxk1Ia/fiFGixKjQCJnDCgUfWnMH96I2RUh7nv5/hzHL
bJelfT6R3wgeoUMeDxUmtoDiD+LtVAvp2ACmWortXJaO9038Gef/9humZmsNnjrgA/UEGvHvRUxO
PiHMFu2QShcFQdntcBv0wMPYKnUFo2k/n15s1yi/h4U7gZq3Si2c2vCbAXOAZOyLahLkn8prJTFM
hl1I7iUuOostqGnz2e6hMP4qGkUwpEvPMM/Zz7EU2u98iM1NUMVuDRBjvzSHRrevX6csiGpQbEAI
9WHlW/uuZlog/RPll9izm5LohlImDwngdn8XFydOT+e6kGMh6QezbW7k6Qvy+vmb4oQOyw+tW5R2
CT6Amw26DvznTILgr9EZQVG84Rcskch9TmmViyAdDulXsax1axedIZQq+iWTNMq8ozquFimC3jN9
sHEx3RoWyZ2+wRXyij+7AJwAxjZZT4PINntnklvIuCIl96vYP3M1YTEmI6EeT05GI/HakTpDlriE
KskCgPfSwUGO2+ohx2GUQg98AJkyzEljcNfM+e5pvCfmFAGxt7hE6oykWxsp3ij7T7q1tlg9ZO/u
4f5lBoHyWvwWDLukHrxjHAvLc4hvxeChx5RiutJP2wum10BOHubtebKn2YbhNvXZsWQPU4G1Wjbp
XOhDQxU1jXXraz+M3cXTsvSeSPaDkYrPaQVKaVSqJY+Q8UtrIt1L1lGKYgUzqww8Kp2fgIB2bugC
93+ap2EjoqjuWG/GmuO2X4ZBdagaTXPsfjOZi4h8zmLSV7AgovC1G2a6OYZ5oDqKP2xVrZMLtJJs
UNYrGMCnosHXcUcnF6QnwNHB+jTVsY0AQURt5WivYjNseBK67U9l0vj4DSoz00HXQ5hYE9XQyRTH
erwxWx43PNFQvJvcv0Hm1BFpJbqP1yY5mXs83pJK6XvC+U4LOa0kVjYHxLX9Q3PuGCpm0UK7PKT4
ZKF+63SQVKR24+uK5/iOgmp+LKWirk8V1zIh/jP4MryoCEBSLMD1kT+xGM+YOnUxA0nga3zXFo5g
XEmsKNnOo/QqYsIRzbd/BDlR6I87SCLv4UUPNdLek42+VtqgNqM1MYw9u7EwrWJ8YNM63mkl1OFv
2UXW4iEIaW8T6cal8wNtQ0exdQGzHAMYyxxRHOLNDYBMr2GVLWqp+Q9t7UgqdqaskIK0vf0B+gBf
Wec0+9VKWG5ZXO/xbU8hgLuBVTX6eLWgQNV/o+d4wFa2gAHn90ywI83Z1OsyoCskFBRxh5vnp+3P
3Kp0wmujN6GvFrONkFp4mLaSLK2Q1z2QSDbpYbHjQxlzyzF1WsVU4bJ2jXlop/g117HiYsZ5KjE2
3Ki00cpYlePoSNNITPCrz+O8Zt03q6md3L/m2tHfDnf01FkUhG7b3lKvlKJKxV0C4wAUj77Hp0Wg
F5hvSLVWZuf4QT5jlYR68Ai4KJxP2CKth9UfntxWi8uKPcIKOpP7SQqprU1B9LD4msDQQxrzuKnf
Go7OlSzxXZ3DN0iy+xrX69pwcCiUqBNxrInMmR52eTbEJFzZcJgXSInPU1xV1EvI1lQH9XG+t4Z8
lxQXVCDkNM8BEyqGl8TYI79PYSAUmi1fOtvCKkbfkYSF5dOSelkVQWUQhkbH6dgLc0nrJoS5fPtB
tr9sX7gf+t/o9Cng1gNHP5x7wMEJ6cKmV8ORDQbIO2h5z4HZP6SFZ1cNN+xORx1yjIfgB/unr7CX
EGj0GIqcV8Ru4YF38vWqKZGxCiWR5ip+zG6cjn5UnCAZr7qsTXYLP/XVz03CoV7qkbgkvbcPDKe9
9x9ZbnHldXg8ST6yeC3xBG/REr5dw5XXd6N0v/jaCkuWkfDsYwmygZyXlIY30KgcwHCGr7Ywjstw
WyqrOBh6giutZ6YsWNqT2+mBsaAJ2Nb4sUsP0ngxPbNbq27i50PAipT6zTuL+/Ram9crv1rEoZJt
9kGW7m4RU7VDrToNpoJnqR50ZqIyzuaBUdlpRQ8QgR78BrTLy9vadhAhIxilGZCDthnfDTXBmOl+
UP+aNDK+4XXK/d0Lk7ljdeJjVfcyQIzQYdRCmV3g2od3+AE/k2Zg4We/x9Tv8kWHbfXMeOjl1QZ3
1a7FO4nguADR1Fe5/ONnflwGDjl58BmaEGyTNb+ipGLpMMHc2skblpzd3fHU3jZgFssX4/s6LlfM
qfNRleQMB48ZotugxjnERgqcKsOb/JDHlTudj8q7TzWVUebPL7+P8lql8oto+x5Eha+878S3Ey9u
WttAY32N9se2fBshMKS1r6Zwn8nevqApnQkyq0r1srbGm76ToYfA0BPp42+UgdsfgQQO2uYqbHyZ
AY/3sEv8xHqlbnk8hHbXpfl/u9JyBEIhQ/OO/XMMQhi0lPPC00ZeOdS9w71+1muvy7YZDvoqtc7h
el9PJ4qY6xh4/0am0a+fTC5vAHaH/bAg+hM82eIQf2gnnSybKchtJypGMrmwC4rV22KVWqYL8S66
z0S8ADKUVxpwGeqBYmymoyy9H1kn2Lm/mxsnZIqoLJBvS2P5vYkF/F40T7FqA2kiFKHhvp5EtPbc
5w4VTzlemW1s/4Nf3sEwmfIUZY3xAKOcaHT31pY0aZBEjx1Ylu6/iwT6jla5Iu84xul20kouFcha
osufzVEa4fjILIrh1MK+dcoAgujAoB09mVNcW8lj4XCOdqNWfwzsk6W8tklcpk/OPb+SmVvz2dwD
SR37C060HUlOtyd++cEcregOI8T9hcyS3+xNi/GqBlVP8IKC/zhQmrAY8dssYyByLvF0St+aAvHD
BPpzwEZdbE3buOaknQZxEIN+LvBB1udeihbJEPC+YAZnjmJNb5vB3CpTXQypEM2tmXnp/4bP5IVM
cIo4yGi5l8IDD5t13JrS/v/+CSx+RrFXFI+9KoV19qhZttuqHuf/Kef8CHqqQ2FkxT31rs71tVRb
qWv9Rkhv+tSJfnRoRUNbXZm1KkfQ+kmxYfQBd1qLy5ho6+/8jVMUer9SmW7PurjUrNjlniCbpTrl
6eRbpFVoOMDalnx6udNY9mLgKIDspR0huZbFNLepr6MO7P9VZuEFUbBWg6IgaiPbO6QWiWvl1ijA
MPP3qNFd+qFWB8A44xmZkaFnVU08cysycWE8fZyOX2CR1KoBHZDTvzZb0Nlg65LSS2D0KsUxCMQ8
0N90JwLgVaVphgK7UmZtvbpEt7ge7hzkIBbl8utx+WN3ahSBgnd5epymiJzYfqeb4fR2Dg8WXlwu
EsMT1DHLpqSV5vtCeX27IKeYJ7g7aAL/ERxvsFqnj09s4DHe52+sDMeZS8s41djV+ifJbHsf0lRU
1qINVx85YsaWZmvjVjEz8HoXtHnFg/PWyxmG6sx90YRLGo7thJTheh6zoAAiMSKXN4EZ36gtDx5y
h+xbJqsFLHgeUfE6MxGdJVcif4KUSNUmT2GDG72R73HziPLSzwAJbvcQwm+F8NyLklaLt48D2U3p
wbCx5XuK3TPme/iP0DYmivnQmJvu0HGejUKm2YUZixA1vpXA4s4l8iJ+qF0b+lTWIcAsi/E66zo2
9/n86vzCwOudzAM58KBvUoctTu5ZjlNofsTZznmn0Rm+uiWlEei3cPZNFJbcScnS2TN5QoEQUHRz
KMH3YjGZDQWvR3KaWCSOhkQ5vigPrnSm3H9Ls1zZGj7HuGjeU6bre7EYwvc5+sog+8e2PPVKvXpS
KHktPu+cm8xpMV2NHLJ8dUznqiLbgFVHaKT2mt04ie3Q/uoIWTcpCHNbVos/pBiiEcVyzSyGMsAb
HRAeQGfKlVdAPbjvySBFvnDDl85oZ0R/twwvZ08W+NnQ8Wa8xQSo3eW91uAPbzlCmp5xTmsMby6Y
p6zbL3f6C13enbr0Sc66fOGjOH0siHBG83CP3cjynEHYgaydMJNXmvDgNBVNMZ4i5EvvCUxuEvYQ
1XlXTeDsum6ubXJrtjMtXX86i/YPWtzqsf7T7zaWeOyk2bp0j2EL265D24jiUbX6VSNO2jlwysLq
iGzu5qqWR5OE5h9JNPJaq9wkQqTBVwgpJ7Jb49ZM21L0A89rIvGgGL/jKOG2MWNVutbggL1/XcNC
qj0TE5FT+ZOO6X9MnhKaoF9tHjgwz+rQMDzP89royYmBwM6EtekMuFpKKiaQPJYz1IR3wM3VthOG
GqqCwRRVyeBth5UDdHT2ERFU6H0tVS50OKJnS9DTC9I/wVg96SgFRlaKmxi+cTznZMYgZnOAmc3Z
PFfbVOP1h0T8IrXM7WCfPWNc1Uh307bq/8sCq1U3LcY6uNgcJKviQR4rNtU+/4Fu8MAjtcBVzlFP
ymy1MZ+fAxGlgIuUKvTvZ8mmUvTmUwc0auySQCWM8aOwgmaUvq5iCylSOUGZS/nZQyUjDl+3nzDf
pj+J/uY3zcXifi0W+8ItAAqfT6w3E+zurqYGaqlbrMgYbz4Vx6GoXxfBMQRpAvSiSwd9OWy0fw5r
yvTTlAhqcCCYn+2iogEi/qYpaw/5WufZ3BUH8WnuRi5Z6u/InnCfpi6w6yfOX/2xOaf5JLbfAPc+
6HTviggzfDSau42TJxS2XtE1IBqTRkBSlNjqwUu16qY57mAF0rRLsUzJzoHidCikY6DBcOEhLjCF
a5CiEdHXTsX7N+LbcnSUo3Un4DPMVBy002SQ65fbrUvCAqTlxENQC9E0XUezbflpInia6vxBUwHI
WLdGxI4lShUq0liH+9sQlJEDakFxE0F0xTEWWim8PQrXlsQmgqdQ2WhAoTl3L1/MYc6TXOx0X8xy
wTA6wWq2B952WW4rB31P8RVDooSbT5cqzIxykUb0GXJ1y+ADdAJiETPc1lBe79XLa7k+ZkZEZ72t
4FX6P+TT+ejDKEYo7R0HaSjXRQH3/bRN7DPnP7PKMg7hWsNWs12VhXgg6evhBY0Yi4iOd4dpJ/aw
pffRtO5dlGZoWnc6JA3/XrGhH81EpD0CXl12inOpFxRRDiv78w0J3LAgjesQsaPAmpv2yABP6cYp
h4JUBy7whudVIB4XwNYNni7d5scy8X7+nhlV7bZVwjnpb2C4V2aduDsWV0LrQ1msKUD6kP4aCYwn
xmquWGXYcxjtlxn6e2thOj/4ugwM+tCl40xuGEXjONFs7SPjbxxlaFVDBB3vV3F7M4vO4o+9o4Kn
JFAgk/ESyTM14IajWbTeiMZCWWvK9BY3Tvf/KVRWsDnZL/6UnvV5iyy8u3d/sH4vVF/5bjDQsY9E
LbzmjYUxv874lvTsxbRHJ+Q0zSQC3AOw7opwAVZYDSTsF3SHgvP2Y1vN0tkiI5v45Fu2/zNSTVVU
6ydNH/n1iBe6kt7dlxDQTfPaxer0lyW51UYoTDgMACP1UB71+nL/T3kY+bkKv/86kXcQzleCMKkH
tw/Tt6YaNOYZPVaBCpZSLM7zg68Kbnpgum+lRconYSfRems026yneB7/bDzkGVPnVzDEBRwuY8A3
xqCvNqYtNQYwKy4t7kWpHOaffYtJBh7or+g1WF5b6D/r3CWyT8uDV+CuJYPRH01uY0uH9oThkLea
gBCh47+YBf+9KgnyTlVi4vMVabcPEeAQLCF+mOCm0SR0PyXYV5C0UZKOVbSY8Cr7BesMpo1ZvHz5
j9/HC2XeMOPaDonvZ7RyjmRfbiYjkCGpv2FTW7ugo9jL1YnuXMnfrfsi9ekZOp6koeAGS+MDE6yS
hvdRF6FnSCDst/dEcTvAZsAbGwhUjLKXfY+Oc5wpO4BvyGiTa+Q8PGTd8NMb8E4Mc2bnPjv0sgBj
5K/rkSJM+96bPO1BqKR8joIkTEFEjSoar2s3OW9bRy5jCDiuCIWSGCgUTXjeI1C9uZmYbNaOZIDS
umkDQxSVG5ee0kGsYdynjIhND6A+d0W4IwBPeaWHD3WhBqiDO1mY0G/dtdfrXPgrfy6G2s+GaPaZ
KOWQYjDhK7WwwXbRsojqZDm7FyhG1ZyNilevElEFeIZN3YyNQWCjFvlSWnp1nH49TGmI8R3u5bwp
+etVXWRTaN6shSfeWxmSN5LSDTxXTfYYULLJtzGqi1Cd+nbsJqYAiaSGFPCuA/5vTDEnk0wpdd8N
uTxI6sB9cQ+a8PhhFFhzen3NhLjIElGxoJidNA621YnYphf39xEY6jI49PY4Xj6AGbYfmFLWq2Zv
5dy4ayaZKkb+bs7qycyJveo9F0aDRMUVnA35PO5o5slUbmf6z1xAimdSjmFS3YbNpxrJcq4tWT8v
AW7ds0I8/ipnNLxU+UM4JDnjZCWVS+mKQhpa1dCPacvrcqrwkjXFl8WsYjYBNjMknzUalzOwPvjD
Ad1MOSDe6weFzpJPwHNZc+zaHR3nF2EX7Ol9x8fm5y4DeclauAIE1Gou8wGprtalu+Ro7UZO03Ef
P2CbFQiliiXQK4H8h0wjDllXU6gqLJBNuLq24RK41fMZWEbd+pZVtQvwCMDC42rgLftNA127bm5J
Aty9CUSaXEHE4kAg5dHDFxYzzAMjXYXYenTF5gZXIya3zcR9Msrd8hv+x5fx7BKc0dEY5sQBBZcT
4SkTiqwGZvJVltPDQ9ZQhVNCSRYi5fqPqhJeVlfT7dfthhZ0AFkXXfLE1KISCs+fBRGXnMDvOycu
erS38RfItGDfbQIrVFr/HgA3q0YPkEpy9sdUvdXkhwNOweV69geJTC9YFYQVAS0Fvb2jH1ZNK2Kp
d0XXMMcH9mvHD6cmTPYNaWHT3qiA5qBfomTcWocmed6pRHeyWD72S2MVyh+7wIGnf1P4/wYDCdAq
m4B93ENZ58b65vy8V5ufh6G3EyyQvR7pFZ0yGA0ct9fXTWxw4HWThstg4bvdu+ntgejOEbTdAzM0
OidTX6bqLpxG0ZM8xnPVgupbJ+3EA4hs4Lm8lGxr+o5GFAPva8EYheNmne6W3Trl+DWWr+sHDTka
WUG2a0Ul9/2v30spJHin8TpvyNBwmS3b23vNjSocsodzvUc0THNv34a/H95Lb+29d03UpyD42d9A
MIE8HBVaa2CUBunpdAe47qVQI3KVNPT55Cp4TRbshcLNZEEWk9kVXB0p+8OJwqFUOut031eBww5k
aWQHNmFBvZTtR18OpOuHiz4S822aUsk+7hanSHpFK1oRzREEcU8CRxHYe3Z5lvAb+bFIXiU9aDcy
WhLyW/4Q06cJT8uOOx5RYulus3v/1IvcR8SC9cyt5sNestWYmmBjtYxyIEv+aEK7CTblsdd0Qszk
xvJcYiTXx1Tn3kRKkTlG2rbmd0Fl1yaVNLEqdNA6j0JnAYBoVh+SAyJu65LxDLmrTglCT8K2pWzY
xxIr86jOl8q+khRAT02PY1HW7d4IIetGrljUG4T2y/TQWTup10G/wjVf2XeAeWT9aKQ+SSV5V13V
ygvosIySRoTHZtpFFV/e00u7CGhmm1vcUmeZMcY8AEcJtYHTmn7NTAhwnZPb4ebdysYc0i9tzFvY
W8lRL4kbOvZQW2RQLZms1evFVMcYWtlSiIfXaFHcJitaXBg5l/254Epeky7NK21GWs05Z/KY8vBH
KPuq/DQ+bGFDLunm3urBnlSIR+gksb7QllyaZPukN9BEWtGOY2a/g9XnlS12PYjRkc2nKN9uOF/5
knV3FeCkU/Z6kWMSVPPL+w2Tm1X2z//1LcK0AtCBphBXCXTNz9C0Omqa+ZXuCqm3S7Kgmp1bclPI
aJCRCqWQJWX4S6bv+6Gr8Kk5pl+NoCmdFv9ge+TDk2QBdOmiGXplWGu2KZHdz3KVJ+Cta3JGto/9
NfTkDPs4J7cizXRJP5UyvK2GVmOMu4lZbRc0TPfkoK/g+VdBN76rW/9GVtobZIaJUBydvb4gMxy6
ZEfbuNEfFemFXmpGAV59nS5Dxy2p6X0eRUuAd1qJuaJkkOa4C/FG55dwAD6av/FoEr87/hTYF1eG
JIurSDwsmWGE6f+6nJMrMxwxhErvv1AB3uLxxGbpIl7WhA3KDG44itUqFJLthauaVIIEvHcCv1io
B17anGsQ7wf7r5NIDvQ3wi4czDeYCUJmIGzNT0Mbzl/bbsR9t2Zxd9Ol+c5rJK+5jzZ/MtZAvlLZ
pUOSb6ArLJi37hEHzDqZuNrlia1LttRKX+Q8afyxtEta9/fcTrtdSZ5ttWEO1yxKxOpOtbNkFqBy
P6uGv//Nc/KRExsB7epD4Z4Kj6g08z3+YIt0M4wv5IJ45Rl5KmEM/WLqrEyVGA0w54tZUXsGX1H+
vxyAVtFNPEDzTzycJkBZ+xYsdinpc+EZORQ0Utw3VN1fNbG13xO9qZ5+rAIhMIZgz0Ti7zQYKDEf
DJwe3aSIc2CIed8/4/IaijkRMAKR0xjnV3Lv/pO8v/r9Yn4aDpBOqlNER9g8YnI/OiYI4I4LOoNK
YVDAnWiKFoRX30knvTZn2pvWCjSwEkhFXvgBNC+pyw1pcP3U3wpm5XUdYoBy5oMDf4sdeZHZGBAX
04T/1d5KO26f0vtzqR6M9cURa3U+Bh1aUxrppl/UhQxG4eIiLd30KdvyElI9odft2kn/QvfPJWHz
p+Cy+y3Fi/gPqv08LBoKKAkgh3jTTvqlSJpJBxC0jz+TJDDsG5hsytuYh2fvmITaxi6ie6ogq10P
4381g+aSrO/rSnWTSjTYmGTR3Q+aoI5krQDSo8cH0tugpHxsrVA2i7/KpQBnWkANXE1DFzsIFELo
lOSXUHVpCzg8NFi2ahODxYSYAzGO5mscZ20wSLevA2WH3OGXtmvRktEYTLliAR5Bvog/WrcvPAH/
Cy3Fm3VVtskmD6xRvls/+QEhh0YGTdkOo4F8k260DPjiXQqbqs4wKQOHhlLHjo/UN4hceHRFlyDb
Pae/GCHdClmCG67krzOgPOZKgr0fiIejZ3KW0qG7ipW3XrbQGOltVm+VussoyQ1qWN/wLoQ6wHdS
bdY9hFmeLYy20lEHWI8gr80oW8UhLioen280YNV8E2t9abb7NUCj0JKYF/qQugv1+NvElEHvCqTW
AnvmI6qaKtA+8hFevv6vIbYql5yjIwM2GG6BtAVw8QULS4NswGcRObmRj2lANHuGXcdPXEM5YqV1
hU2qJLsB1hO6LcvPC/3piqPR5XIbc8M0e7QhPJnATb92DP3aNn74v0E0UaISkgE00wf8hX7NmjoK
ZozNFWMZPTCRZg0RVPt0hLAlnmtSL+bnWzpPzCeFEv/8xrsIOtZXyNSR7apkNaY/tF8WBFMDQkVs
aDJtnb0g7QKkw0QerT+ICRrvApnJd9mv1RfetJYS2+ahXo+z+uU/oA/GvURzybCdKhP5Y4qGNqL3
7JwEMSYFzwk1xc5PYsiHv3aVhONJDbhfhYzYF9xAPLaWs239R/VNHWQlmZ0zlnEyp2dCbvAXPWJu
p+cmigT0mOzXGgrPUXbzuHaUHuwvK21qrGu/vn8OEoYDzXRyYaHP45s3mUCQifVstVpsfuLf1+Kd
XwB8KZ+yBQ1sFKcTwJtxqOPuAc6aVvMM23SiKr3Pqdb3Bi05ErNMKeSee2RVxJLtQ28VzEO5lut3
Yo4Iz+uLkngeBSAha4e7FXcgtFtZbgvwkt52ALYRvPNCC+V4VTiF4gkh0nsN8mVc02amtgKIgMc1
L79HauXV9RbeZT+OVCde6yRYa4HeaZ9y1BIvNUDEe8qzDanXYgoMnfwOWo6B2mEzDI4Q/C1KMaVu
DW/Rf5a5wEiVfNpllYPXaoZXS2yj7rzfm/bPZ9NxOsowWroxLESCLNBWz6RIOktFtN9aH7Qe4hqG
pLjZ0d++V9M98sGNcp5WLvvAM9G0+3hjuulri1Mb8P++atzcbnEu2UEhGkgTijCHkSCR656pqYWR
U+IJU4/j4YClqOE8dO0fJseqn53Aeh49qPcHjcqvzR9WYbH1X+EQJgWTtNiXquMYY7qbu4VTrq+s
d4o67oxHjBTatfxw6qowtzWkXIakov+ZhfDX0R2Uhl5ixiqcdN+ZfFuWbhLR2rgJr7DalQhYDvD1
00MGtBs/K/zz2Iw6ebixZGEq6a9SDSq4PDISvqwkC1brCcg+oaLe0h1Oy0JlCNGQLwhUAOvfUJaf
OjKaAe8rj6jkukKaS4FBJk0++hgWCVTYl1ST2hmaowXy0UCBP9k/yekDOqUcQ+K+73RdD66R2Twc
t714gJVD8xyMILDAxiahLo2w+pxWdBsDpmWSLYPG02TgMjHZl/kRnjCtLvEXBLJrEGcn67BK91Ci
vNsHcqfRvhyc/VeY9IbEGJxZ7RXRXp3dwwGrESqdENJAAMdjtkTs9SgCi1PnivjjTBZqjgwhAGtN
wb+kZyio7xu+ixk2KWwtSj01uBnJFfv5sg/Rcjx9QEb4+khFdTN0x1l4j3k6zmsspQ3eyM85u96w
fsed3iw0zQKbN7/9RC7ngA8g7hbkCmFBzPuTgIGWZX9+LvOnjb+karHQCJ7UWSZJ7dxEEVxqvS0q
lhQoooCzpGGRa/GOMTXk3Ev3UwCMEGBQrGP/OULsxg8YZK1hbMKsjohVwhifQ29BYmt7pWzK+5Yu
8zAf9gtGZIMo6TLaLiyGCFkonJE95ShMURah+4dNDbjkGSg+6MI7IQdJagN1Gb2cJUTP8wJLEZ+n
98ktzTRrCGdqDbWZXRAd8uZTdvCJdAs8sm9WnqoPgkJSCAYJqbpuAllh4NO0wRIMxR/j22mTwc4Q
Qg3v8cpuxM9A1xN9Sje2Jm2D9i6vB9MvPL+8DeGz3LSLNgw8RgVjyouaDOoLHMm5o8KgOMLW5x4u
eYkBPgZhxUsLEap3mNEIPSDVxujArVnEtZ4aDPbdl5CnYpOJ6u83RXcN2NWc6C7be0GqGP4K4o8j
kTAXko9OcXeuSCXJrzjL2VNxu3kFrES1OIl61FCu5wqJbhmiyVL0bLqGp7Qi65gmiV3YiWBx8hX6
jmaSsmznKpybQauxAx4ZCEloULYKyKvfz/bbomug517ePoA4V+TqS87i6+6pS1j+WJi65ZTIiufC
UGOw0u2SPkzGLL0D/qJDLXPGjiBDr0JjCgWUQcjJQ/G1NWYObiQcO4YmVH0bQklELgnqUN/PI+SL
ARREh7qma4xb/WWO7UWin66+x0DwJyrJibG/gE1yen3TBgjUESm8JnzGLQGC5h9PbPSy1W0rENc0
oneZGBFrevneMFYMgLhr7oqZHHl5KA5yZrY1RP9JjNblBVZ9G75UIbzGbElIWXU432C3K0Z9HEHt
IUS5wFNo4AxtZvm7rGa72bHNJRAmVFC3Zb4DyNWIupU2Q52qoVmd+9dmgyODS9QWVdfIFCrTMHdc
0Dw8BJIxwpEj36gqpM4V6gnt8RXsl2ceQOW3rP5V+TPt3xZKLnKr2OW0QrGixnQdLk4+fYyUy9eh
wV0h1mUo8VV4nqzDYP5ux/YDhP2TkDCqWmD/3c6cYUzoSjGGQsIsi/vkSluJtSq4mihQaxaBOG2j
ShM27Y7e3Bfjjjnj4FUWevZ4kKjPbQwRclQZ4lJtjUxzs6prfBLjpCTi7rwQecVgA16Z+edUqUCA
8tfVv+sTkio6ywWirKsSaq7nqRPOVVeJaH5VmxmKnwtWkxeFwmOb7xLhdodlPo1Jk76bur1Bvvtx
G3dp3e/MyUrM+mxuM7zbCPBX7na0VO45qosUCNFj47lh3UXHNPbwraTxBgcuDOC16vyNGlz8+02a
sZeWixvxmJVogxORG2kg+OkeCvNSH7QUPmo7IRgyl6f0r6upgFF0HFqzdR28izFBxYb9tIViRHH/
SQjsaNhHtiD0c59hpvF1+Gf2ntD2jjgCSlrWxf8d6EVxQuTWEsoVPo6sme8WWIvL8qRhgWTlykVj
GjS0ZvLhkG+o++j5XeK5qDE0QbfzGwxj5oZ8qRup2BjLQs+/kaCZA9Y2wa7KIwPBQAPXtudueR0i
8WKjs6H4j+ifYsT+arMJYqGaonKOsSBL4slD3pmSrotkiQvZ1O4nghZb88qM+Yqlh0xlPUBED9P2
98fozkqaPhZBZIz9ML2jNdktBAPA9gD4WY1yGX0/C6lzK0owSz0BEb+DuzePofLE0FqWzGWZnIbm
rmzpfb9st5U5vn/qTAX5Ius0T0C3UCnXw7g+z/HOa5omT5kaqIwObEmYUjBQ8BK94iU4BIClBZ3b
XSH8FlVRDnOrO12hmMzQcslbqSn9egfBJVAITYo1t4zJ3VvZvc0gcpMBcn8X4YMy3+vwuIPRxr+r
OLyGRHf5gtf5P0ZEPw2Gp8OiU2pWKFW2okRZge18zeb4vH0SHqqGn4Z9lYFe4fM0tHTP6qLEfJzU
DZhRQ3JEyaINdjogyqcvCL44aMQ02lwhPvNY3ESZxJ7mvwlPElivJ0NxrZdiVbAOXRQ0rqoPsDrC
QYAAETwZ9MMl06Hah73l516rXM8RJEUqQeF25zmtfzM90a6BENeWat69JtC6T+r2V8crNeyGuOuP
Bml0pcT+DScBhtm77ExcOonBD46vuBAM9cL0a2gBg/PUETOjRyVrkFGZNzKZlEz15yLcoG0SKjkX
gWLTyiS9xrhyHw5rDIFZYptK24USYBMtfeF1SDDRFvTXITodRfLlJD2JAjW0QRw+ZYTxHFNayIUb
QU9+M1dafkvXt29msGdgLfGIUCA6zPMS7OvCb3KBXxWNBoZqGezuUprrlQpxybf6y/YxAbbPiZUK
vujIewVQwkj01PzJYGx7bhzYqP2dWK8e1TXj3HfQOYP2sYCVN+GmqbmGtPQQchVzwIF3QKgJHPq1
+RSRYayE+t3N4bkCgMzbUugTt3sMQszEon9zYdbYtAOiCAr6FqspRYMxSHOkPpcPI6yMoFcAyJYL
Vv0teY6qt5voDc1TAZj9xonmLltKz45kFePEzibBQdbSEUnT0qeLQp3WJcAU2lbyXYKvJNCXddJ4
VDG946wRfUvoIC16TAEl9XL8+fuKiXe/o8eLHlH3jDMdawiZmwhXdcODxrHlJ4hjxGNsJCdm+UZ9
GanOyv9zanfy0kR8UNK8abejzmKbk9gKfVPrRzcDmJK58U4cg6psyv7R1Q+MjjyL//6udDE7uXcj
udFeA3St1h7W6McYvZ6OTk+bwqg1JTYkW/Dl7E2Qzv0e8ue9enGxO6YvAuMOBYg8rwsn1LR6A8aI
JRWr+yLmSNirZRPUG9qf6rk4btMYsIsvS9+E1YJ4WZCrrvZdLSfPAHNMQdttUnlVgzEhtocp/wGo
nQq+cluNXdmHCtc0WIP2fSaeBVWTOrQlqsBm9yFznRlNalpOdCGtBFg2DjkQUl4z6qEirJpfpXvq
01qsPn1Z8UGgF6QZlsE0AFUDnvjM1rsMuLx/OgHj7aROZN0Wda3hH2HxqrOWh6vx/G/w2hEfeXui
nvwb1zfutDk0nYjVFsmwTi3VveKWsX5zQ6k7aCUtyH5s1V5JR+OAeSx9FgRuFDeKdbmwK4HziULg
gou1iepmOvWDVeXOoRXGCulUrvAXjIQt4EOQOqbqXdgY/YQlZlitSWnFlWw9VKse3tsDWsjGHsZi
z4qHSv/StgGjqbh3PYeZ67v4KpvtOFQ2ME6C6jnjno0z3Ke6QTNR141AwC8Onzv/5Vh8YNRKRPYj
SR8z+EwfOkkTKGxxXB62Ibo7vedPWc2TDAMzDOfH0athK+6ZvP8a5eekY4ahjBJooZF6DLz2SvVD
aAiH4zDwZhO6fKiBx1gFvHCftnM7SH72ZtoJHNdbascRMnlMBQNTgoWVSmXy0Qwnw6pAqGMndLyf
61o1QlT8RI8+TCu0hS+6YslMeMXGYrE/QJWiNT5M3li5tAsS1Gc+PEIkvfI/Y81+mR8kjd3NlN/6
kjquw4K8gSPNcvjsHit8TV5+TLdE4VF68bv652tZh9eXy3zhTlCmdM/kAr2pN+XiX0Vovtd/ZVkn
iXWNqGN2tOSXvi0Mi9W26ui2lKlmZ1oBMo357PTP9mSdso02DpO/C8vWHC47IGjjHBzzjZ+UnK6b
Xs/jjV5Bham/7O2oqMiLAWSMEmMN6plUDwDkRRa1AC8Q1OloXsTrKQXVYmg2J0dyU2PQ+gG3Urgd
0p6ZCIasz0LpG53LO1+4ybJO6A0dPdVA6avDw3jLpwLYPv0mSblSuCpwRDv9i9d4sAiQBJpfzqlo
Z8lyqHZWAmAzSYKIzX+xunLrduY7Skuk0REskOjlngzqA52tEmNo7T/ZtK4VTM5NVvl7GHb/6BOL
TBq0Lby38+QEuSpABeIdtHaNOVgUdHA7mmXxC0R6fKMmJHb7yvrWAHh8Qdg2V1c590Pnf+BwIUf0
33omIQ4K8xXojBo+V4kgYyBVO31e058Ynccu2keC0dnCq/a+UBQcBh+tuQHMTWGkXXCozu+rD8da
tegiBBWnBBRMNSDyXX19DCrIuzXJG0Zk3YbcCr6MdrTOV/CHLLtS/B0PO+j2GMhBcgMh3EMVyPVW
Ndasj4ogCWPjZMJ+I0xFhKDogDYLMQuz6dtXA27YF2yTabhzQa8xqq8qQ+hQUw/B7TId0UsOKucT
OlWj7YdWMSu2IZqE+F61D8r9XeSoP+Al29e777qFwxR41vw+yHA0dok0jBDu1+qG+yQAK+C+CSd7
3u274qia1xT9ZT42X63qBvOVjz7yZ6vKQ7tedA3q5cwdcefkAKcNB5RoE3X5kWqD0yEj6WmYWTmS
WN78nxdrzfLs5/KIdgCAhUAdCW5IMxaz69HeD/NQTLHN9hwaFwE2n90qB9QXcoHARTYtFURaoLia
VBM4XvdvfqPi5g9JYVKkJVO+YywCvrP2BpdhywWwXReLNreu/FlwABjZPdbydZCGvt/ugEymK3d+
of7bxj281f6bzUEzPZULyaFdiTbLEpOywNJ5NcL1IXv4cWmB8YqLtiC7nAwAQM5gQa/otWh8iKe8
HA2pvSyCgbiJVnnODQQrTxXkRJzov++2yR/BsJvYlhkOwtSO/zm+FOBB1x4l1IInMglFxECg9hn3
OPmRLKwCWur5ywN6iBZ0YXAlcrfsipxinf1f6nuWrbL21K7jCGSlb+1egC7mLbheDeaBbPhqin/n
VipCiJdvTomC9fMFRgE1Kl0ckwRZMZGTaPwm3dGhspyzYXQSHR3VYduXpTqPT3ZDXsvo7RQYfWsu
3r2Deb14x3Rt4J8vyQc9axTYuzNAF9i5fk3xAW1wNi50MPi6qeShWnPXZ0dtIk/UEk8StBb9ZDa2
my+cifVEHksjs0TfGrcuv8Di9Tj1TgYOHUTlVoSYnkcY7g1/5IHuCukkgLRyEVFLmHaAFdjMn/ic
viVg4hUwAldftDV+A7UHsPq0jZXRjcmeSuKKSB++V811eSDiv+1azPuLf5WwqNEUekSun6SQIwKq
dDQ6w+r0RlJJwqBqwuIlxSqA8q0xSfMzCBKCtjxE6YUkY674scJ8vY3VQ5dTxVPtQoNxS2dcLVJX
jPm60XcA+Ps1fjPxGvJxyjW0fBihzLZGmp/RgZ+mXaK0MBjh2q+PEoEqtk1qFAhw7kyIaDkaFs0C
OKyiXAYl9AsX+MQB3mkQ+ysYmDzFZ5c/NA/2TrkpNN5PbalNLb3t21eBIftbgy3Xk9YThsqs3tmL
uI6rVKTsKnKFjrPPwtQ3J61c/5sOan8ymb6KJxsF/EzyZDHGZWK8TDD8V8NAbN+wZdDR4iRWR7RW
qXb40Vfz6Iz3WY5MQF2+JMTWJ1rOqLkYJqGPD9cN0f/MmA9kiMFEPG12EERjNRQ5wsmsh5JNDGAz
kzFBsSuudaS73tYaSwH6SpfvObxNkw9C3EkI5AQtPxJYqULh6DefL9O9V7zW8mzqcmSJsRdDCgey
K7N/+P83nAakZAsKwLD90dRW/TI8KxuC38qFBT9VoEDtrA4kKh+JY2z354+q3/xXjUzifWpOh5Z1
To/dm+1z122qsaacVyfiFmtEC/DzppNi5NpbhpSbaTHau6t9JFA+AatjgliSmL9+hsFLnec2AhbB
572kh4xcAE/AjU4TwYBQgJk0ddc1rsrcl1QMirUus5MZaK/pwACOO6y1kWlCcx5IE2S4Rc/uZVuR
7mY6buB/4J+Sy+WYenX3O0PGlKAbcjILqzNd9eCDwEglQ3q4Jd0dsepzhK+m9/Ww8+r4Oz9ruGqf
DHMGRm+xSZMDOgMVhH/9gXyrVnMspf1VnDDSABw8MIqZ29+2veyMxY6S2cqGADp6bqLsCTvrpMFa
LTiJRPRqP0B78RGVsLFjbfkDu9tXO+VTR6IqausAs67/sC2OYpezMYhJaHGj6KKMx0r0ulGpgiMm
QEaTLaJC0uS3e11UQXxV4LsCEJe6hHhkyTiqDAesT592y7c4xa5E7j+zUk4KsBT5vqrJY6IL4RrG
gJGr2FathnbSVwc+aXLXOkaA3C/ovE4+/mAKL0q6QVxHBiAXMwEvov/Ll/r+uMCTpRhyYphi5ItB
JY1+QyIR2kpIY+eP/0BHdLSRL/x3wNifRuHvVIj8aE43GHZzakg55WJqRhLyXffeFi+4rXu7N702
NYkxqtEehtBatP+1cX7Q1zCrAvy6nUAZlwonT0pb7p2xNpTP0sweQqhRNi3AFtbjtTdJBOk1GHM8
OQxPaj8QWl0IQ+Lp1UsEn9GI1xxJXNFVXIdp+9zUOOA8LiHqYKuDEbKzByGJtNcT7DnexaOupP1T
SuZCUV388nyUPCi7ebKD9h3ORuICwFElZzmshwoXTZMt8dcKYupPKbP/hly0VM2f54xZyJJSLSst
+KNp8rtIWUQ4IgyDLtE5pVdMpA8aR0mHR3IIM0YT+jPAgSLh6s7jRCN327vklJZWjlstJ0RraTIc
L1FVy34dKyhjIO7XxutOzJX++1Q7R38EBDGugZEeGhkcrRuoROlqMMGDmr0Ife/SRddDawMmYOmK
uWRJZ3H3zj8nNcRbPXtuvx0IQ7P4FqhfM331AK1Iy4irEKTUdOdvcYBXoZCHVktZqxOAx9EWbXSI
nFuyaPgNtIStcjudDI0yUnOT/VCtXB4teMpG22RzEE/9zSYD+HsXtU4VSpPWrBuhMYBeg1p6n4Ki
e5K9AKFbwFj/DpjnLncVb5fPPQNVUPTVtiNZ1L2aFk3+ELapWl6wKJvn1/GoJGszAngdUhXL7yVr
JPLLpvlue8HM7tfJiKlRzqB6yGHE4cgUsDB/uoePnRLSvjdMUwJZGn1UZPiP8FfqEps3gMRLBrBR
HA8ZfuZYp/fkGmKrHBcT2gqelX0nDh+3yP8Vl7QIFBb1bGyThLUssVysgQB0i0G+o/Mu6bRvYpEf
DHErBxOhs7GPlMLX5O2VGGfZ077qXsSRBtDZcDuPhCpUbo6vCtwv/MkTfDm8Bb1jBAqw8gVvrNIR
pfQdHRshoFTNzF7n+XeqYFwMka0YG5ZhsjRmAL+isJufKspxc0fo6MJCokAHULfRRPbeqDg6gnzA
CFu2rStfCdRsz4vHf2E3BDWt3p3/httY0gE+51FFjGvpZsMDkSfirGXwgKrGOj8E1Y+EcjnaTe17
Hxp211RFPPFRKle1oizGYpvv9k4Ycj2jAo/vIVdm0hnKvYGXlZVh9XXGYweeXi7CWFROPfaJ5Lr7
x230UQG0osA6kDzUz/pWW0v27+NBAIecuFXrXkVh6aH4Ve6PoxcBS0IQmOdS+PN9Sa060MMjNyaD
thXYB4ScrGSnjBQ1OMPFEhrnMOtsDlYIkFdJgxtqGXZl5gKSxQtKRzAMenSbOviQwWUSZx6xTEr9
DXHFa7xrLV0OyMQO2Yv8ScHICidaJq9sJR2Ma5cbJKhKONURrQI39XPoDw/z3h+ZLI07ETT3EBhg
qGKxytFwNKGJnGpbVh0iBewAybGORBpm25IX6uSHPOZXhxJTV85scCmn8GlPpGOsaIFvFJcj0k+z
EJHYA4vSZ+2SIhr8QFrMwBDu2VBsYU3sdiHzVrEKa7P0eXeBFHVvgvIhchJCa0tqABJjWrpnco/L
yjTUsGOh5YXu3F00+de62gTFB+j5/ZdYjhHYt0Q6Bu1N6aBL6vylzTt6JQZqBFHBKLzz/Zjo/PT4
6I/ALe12dzqj1OGkOrVaAcT9cz3Dr5FHfucW5gT/3bcqpGHqwkdfPuYtHoZddMXzoqPX4sjep0gW
7P0Ztvlp7nnjHMHMys/01bQod+SHD5aZHWBIVKP46N/myU9n5LUHJSGdW1kFtBxAJwL1Clsam/vl
mRwAT1j4BuBVuzzwybEmNAb8cgzRL7Nb3+phFOrNOYG8Ui/ixGDgbiEnfz70CkYcvp4y9Eo95ne3
+3f7OHOWVXIz7wPg5xA+HS/3K6oZWCvRZeC0rRHVfNnyX/biqKoiet7OuF03f001sL4W0UvrKzWb
tYA9DdrbJaOJOUu1rnKyeixoKebueGSGcdLqu7VHYUvBBQgdLO1NgzJ+wTJFs2QQf1uL0rH/Qeit
F/Qad+nLuxkNR/FBdDPr+9q6HHKziK5HdEfpKHq3uWsZfVjC2WDAWX3qhuBlPahiPn6Ujf4ihnOX
uWjm9VOvcXMdSoTNBn4Mlo44cf+B3DxcSEra8DCZRHniYDEu2ZTnS8nF57Vi/ghyOubxY7QB8D8q
+pHg7mSPYUgNiIYh591IQfK99a8QLoWtlVd0/k1kp46L8YBal/R6wxNtl8TqLoC5zG6MrNNxkil4
YYPkMbCmaZieR/rL6fgdgbIzo6y1m8vJ3aNG2jTaJmztta85RCS+rdRUN/wjN9B1LlbnU/rcfesH
LcMaqd1G9/CpC494ztYu5AlMg+WBE42qjGrAyLvtgj5Gsevygp2P7be+t+ukyQPr6F5oZkUabTq5
/2aDq9cHyMDY9gneJKE12ZOGU5/BGMNrO1FutgHbm0Oo/csL863qqLcsZW83v2Qc+W9CVxrQIw1A
5fymC514ebdD9hh7oU87soKi4p5AYOsQO9ybKAUFRrq9FsE53vbcuOiHU9ScNeHxVbC4/LnKfgCr
GLcooYj2J/9xee+nsnKd2KiIYr5L9X6JOvQN2rmG210Q2neaGnDLNC9bqy2Y9dh07cgnQL2c9mFp
UUc8/B8RMqAfbDlk1XVwS/VmxtWb4rEdoX1feJvfa98KPF9XSLDhePnIvEpACYZJpdIM1oIevamj
cU1xwQlTL8nPFkkSLiAuQp8Xs17KZcHjSeiAsseVAKS9nARjbwBBKh/pHp1C9LDb6zrVInescGkN
d/qjiBS5LE0uts6l8NeHZGGya4Pp+SGvTuIRlbbSBgE1sXBKLxjBRzl/DIhNQL3It6DMJ1Bf6X2Z
opcucm/fO6rdj+3mK0kTnaxEmkMsXsCdaeLgvLXLhU+2wq+BUDt/tSkFPgNtKh1R+Ct2IV7U4THF
Q8DkA/ZWKCA7QO2LVqNPco/UMkKVe1j/xzNMC8frVmSKwnIpHSe119Ys0o0cXEem7kvEKhO/QWAX
K0uh+W8gkTIyFg1L7zll671LqmMPizy7tOBZbqEjTcxQzJuMb8KLWdpGoyEo3D0PphXcfsEuQovl
dIc2NbsADyBJaIqJ0/cKDj3hK3aGS0iSS3WhdH2NsPnVDCzHzoSa6Ag4Q8ZQvxsejR4JumDeIPoB
CeS/zPKxE1AyIHFKL2KJsg3woBEGP/y6m37Agi9KHj1p/SodeVpPYgYgOf9uDWIkQeH1Sqb1auJm
LEoSLGUl/AYPyAS7eygGnRm+R7VMHNyPd0Se7FrGFfffQOS6n73abR9QxtqmjRBqBMOGselhXqdq
4uWpvI6zRAw70N8Sd/MEmhfkDLNnX/3D2qnmPAaNtQVtAyQKkjZRVITqPX/GiYgosyzJcPktFXj4
+Yyo5gmcnH5saROz2/ne5Pw2GDoJCWskpxOl8xIKuvDC+v5fyjtdvWYYrrQJ856IrNiMAo3sf6ng
bt7VKNvCo7X8LbLaKGSgiMXYkgqnpTRMHLEkBpxsHsQZJat40sD2drhwtJoObUDlvhTUkW8ubbuM
2BTtd21pRIQgCLt0CwJyQhlDor+vOCx7M0FT0phDZcZY9td+teikEpyGvZWDCS5HkuSoHRZQoWxr
rwIkfrLNzxZYz9IW9uU/T3Q/3+eWO2Jn1068LhSg9SbjW6dusTMZH/C4iThF3zReZqNtD4gjgwkJ
wilW0R1dWT8jpG9H58OcXaisHvG3eqhkrEyVNP0ntIfkF1snSlM97fTPn0x2eX/xJcNEidiEhANl
eXNtlZXG08AeHc9LCLvqWcJVWRutDeCcZ31A1o4IDt3VfIBtAMblit0N8Hzvnspe7CgfVNtfm+1P
qpCxp20Xy13KICbBldDOwnx3LwsbSW/DZlgiVBlXbsflhp0nWRbSpZGUr4VFG+hRfR07gsLii05c
no5PykACB3j9CeTx+Bm49Fm39xRGZcqx91PWBE/vKzEUvUYGBBqBM9ISfTXUnQuR3hp4oB8hwcKV
LNeFX8md47KYBq/Ag0m2F3hZaSfWbJr3Ugm5gnKwua7ZIBo9ZVN1a2m0VxOeTK3+u/Sei7V1sXXP
OWC/Da3RSfraY7F3cQTwJcrEG1yuVhQ8u/FaP3oVheqAs1/93ZnPPAxzp+ZrtO8pKz+gIKahWA4F
d+GiPm9caN+ytc4AcroAvRnPt0fOFl69GgCHV7EdwgWUwTl0JLSetXU726ac1sFfkfAw2EVIwsGF
IdkVDA7cQm17F4Tk5TZCPijugkpAYkk6YYai/OkPf/3mP1jOkqLcdMfV0duVf+wtuYvRPDmzOSNK
OHqqtoJfNTSNVIO0V23RzCpmOs/kqqQ1KqrIEc3cUkBrcD9M/BZPr4nFfSncZP0AP13z+AdzwNi/
fQRrvj/pA7QUsZXjeoIHkR2nlALy4oTM6L0EKJ3f987RCuukkLkF6MxEZFizUQcIe+twBJERofXd
2CNdM/QQQvR9uz7N0GUBTGtUpwIGLy7G5GI2NI3vhldFaDl6eqDpFTMjJVy4N6Rza8CCl7QbJKQ5
8oIxGrLdP6nKzyVUz4SKF7Z1ru7OTuLISBxXuyA1nKg/wbg0Jw5styGx2JAE/S4MdpRUzkI49LIX
7K+YaXqDY0ddgrcvaJVpOG68024WOli68JyVyQteTsKr1IGgTCNAuH8Fjf2uWS/NfRNm/de1Mkp2
j2NvHm5B/BHyaYFugXpXOCl3tE+W/7CRFcjSwCuzILsk97tnceaP+JiV+61AhApiZbZu/8j08kjs
4ns+GNL8mTJIsB7QqJmfm1XAzxwqXFsNWUM0WeCVrvpnel2bHi4APet9zDXPJ7J0eHebMtLV1Xia
c3CT87s4QDV0zl5idnVlZvCD/JOWMWDJOxSLm1WKdZiGfzjt9I/Ou3aMy2zgkmVR0x2JbPWyrm9F
xLUF/dJLLt92ntUt/Kn5EoIWrGOFWhoTlnL9Af8S8UQJSQOj4d/bqOhlOUbLpt5E3lCubm3oRK9r
nLV6KtSNrHAt37OuEOqQjfGje/5behAuBWUDheIY0iOTi7A0lhXTiB9Z0QLQgkd7Hk2BVRfYNLB9
s8qYE1Oi+nBh6DxEgWbamFjRhfe64P2CuGE0DyTzqL29AsRy5iOQgZncu+lJQTCSNHGshsnBnVEZ
q7k/c0To+ZcjQ0KEtNImy7DCLNxbPSdfIDUV891v6zi2vR3mjIFH2ZyRufpuqpsPdbY1UgLB30Ky
m04o/R4zto5ts6oDx2IIfddV4uFF/y1pzpdw7X/NqFyeId7w3CvSsyICLqN8woRcXGDxdoam5bXe
sqIin3sjTXwKHI87FGcQGDwCFR6KguPO2ejtjjUBHt+tYHzV/J21/6XrNAJLizmAfROyREbJZ8Ht
6WX9h2azmW1FLspfsk+10fzO4KaKsEbjE5oFj8r/rNxabdvqNxTG0Jce80Y95HpFyMf7KqjRNXox
ORf4iJxT3EtXhjmpxIaGVYTJa8GBsSoc4MpRdPu+hUXKcV7+qpo80f4qSf+9GqKB+bR10WcfrxDm
vT5KQJUvgcELXRIaH2VUqH/ztBKJZzt53BT3rQIIlNGOJmjnX+EFfaSJcbCtY14k4jKT17HD88+F
z0BBl8SvMA+bsblEU5Z1x+f5EQFcHIMYhTq0i9g2OGWQjTArTRV+076k0jOx2xZQd8hIl9iSaCs3
rkkfPLd1fM++9Bf02rfbGLNE2yiajCv14i4gLqmgoPIXEhgaa/Hr1BxwABGG7JLXdrngEMzgIxxJ
oXjsdneT2dmbTFOHy3rfK3Dm4jiZcJJlwhSANHxwp0RPNWA4j/3T7SNd1s7DLJmbrL9QRO2Jsl3C
K+jRdzHg4rY2sVYQJKG+TxWm1cQ0Ln1ELp97+/UG3PlGZUf74Rak23bGE5HgIn3FQYwcBoHsgrgs
/e5nvBlLwWC8Sb7isqsLLNmBbZ6BgAmizL4nyxpIWIJAT714/I6+vjt/ucR4Ham2Aojldg6B+qOl
xG+XAPMCxjwsm8jV5jfs0Hv2eUEzFDrjgbjR2lzc3at/1C+u+3thSvBaiUbajqQJJENWiOJOCRX4
f2MEdHeQ+2rmyneASLzV3ZNBBvCC5LbpFqznHVYrGGRfq87B6RkRZWKQ/U8UlI1Pb26XI61I0lDp
BOV0mzWX54w4a3IDl9EqZZ2liwYJFRqskGjkCs+p8Eib+Muklv8HFubH3D8/CvZ70ekDxBSO0WVc
87bWaOS4BRdL0jPByGMrnorQZ2OG35YxDUXdAUIfumocj2YiMtqM/20qYqMHitp7/ENxelg28QyN
Fo/ClTm3FpXIgZJ7thICToxs7Woi44YxeLTDevqkuXeDQjfAOfKYNGTR/xoYEhwbPhLdbGHWRLeS
5CYpv+TY2UKAGc77YnBOcyMeBWf7JJOdLP1UPxc8Jg2FQW3G/xCsE//RCp8OpGwiMQ6EmqUcnJ7Y
z2axNzTjeCmx1/2unAG3mJ77TySeMTAtYIIIMyOTuCGzLmmsdtkH3Nocq0xzTljtx4STDMzfJLeb
qWj0tPVmKmkXLynqe3hhIX5/WJ/frrp8EAnJN9D83Aw62NxRzwuRbkf1rH/Kl0e1HQCF8Rskz5BU
GY8hxH8hOs0FT0Okm+ZCCllmGuEOrIZKYLc0nPBxPWjAEpwA6LnnKBZdJhLPWcGK2rNhY4PwL9iH
1Gk7UMG8Ew+7JCfztQjQ6gaOCn6TLoufUexeUMnpwQq/l9VfDs5GYDo1Jp9HAqHcKr/PLAkCNFaI
g3tlH1uOVFTgf/lA+XtIOUs8VBcPWKIr0RM/HLEfXAJHXJdO0Tcg8j4d6woev/jSkp3OzTS5fPa/
lSdE+oPdtOGTPH+jaHhypVkIFZhfLd5BACDsDpAVhR6geb+i4Abt1rvn0R+Y/Yiu2owpSFZOrugA
rSTM6LhYKxKzzgaO5FoeEjpJdK7q7Y84lxnQgDWFM1sNu+meJMFrFx49cWjaAuCQEbvWOvaQ1yw9
Rdq6DeACKXgotznuj1xS/QXTslscf5jPyl+JqtLRroiPnW/tQMJko4JpRJ1LFdnHUL+NuF8XyurY
P8HiqtNtGZWfo3XE7nGUEKwFOZfEae4ZYUXwKNmAFCZHlr2WOqHyN+RXeWK5RkahLt7TAFodSLnX
5DX0Y2+YR7Y88f8xjwEiwk8pVJVd9RrCmR0PxdlctScMrGcDsrqdHE8esA2aGM3EsedoSyFHd8UF
B5O0ChYN7tv6uVzzAUhOEtTOPQqLfALp62K7FqmiY9ZF53Vh+E5gtPyA0EWgxrC8616r9QoqjrM/
mHWWCH57p064Kijl8bK9T3n65ZfLF69JOb8v3B8AeYliSBnQDY6KNA7+dTNVn7d8Cm5hnFDVsV2g
3Nk7/2sF4bXgRBtgQPBxDCI2yys/Az31yYkfDdFCoC0+ceVf1KpGyx6Ptf7NxbiW3YM98DInknDB
FfKD0KxcAJKm74VU/hCD04DfbgLriKRXpMU9AqEeeJfis2cYqSoPy/AfNlDzCRHKIby4CirLH6TB
BZwa1MKxDyl2VxKMMgzgL1KY9OwzYaOp4BArEfzX3q86ywyuRQWxDrneUYopfSsRR9hutkH9W+yT
i4xHTtRWR2r0hol7AeXqk/izlcAx/3Ikwk5C/+CfffQN/erGIbf5g2Ngp3yi4fsPnTYWwRNWVqhy
y9A2Wp2zMbz5CXZP6OBOT2BSyfP+o64VbZce1IxRWghDBLIrg9nALNoT7nbwA9aMsPnaX8Tmmtdd
Mn1th3Nh/iF1deNQfLtj+6h/DyoB/X7hRxMhFyP4DsffVrdiJ2SugYC2m3wcwGhR4+3uQw3qsDhF
Y7J4p+GIqPQzz4mg3Kw7z9Co3MwhuAOYCLQIQBXIXRKPdcWu5Qm7u/d/wjVWbGTi93+mlLyLTRW5
feSOvkOzs/H1stOpLa5y7mxKvG/l/cLUilW3n5p2R8BKXuEHXvVMmeF7b9iw9ff1wlpgYERUdeYy
t0vA6I4wtDQaRhQ4UgUvvDbc2fpsGvEE5BDmQBBaXVc4p7C/2eTKnHi/i9PMunYOHfv3RH6jcaoR
SB/l8uYFp7U3qSDnr9C0OW9zttLdhw3aA7ID+VK0FIY4F7imwDjheEPdYBxvB+eQftxyHx0b8mwj
UiF9YpIfcQXl2WSR4QYZiMv3sbOYX7eJEfRRMakLL/s7SkfgM6sKSI/N81t57wp9iNdjosBbHKIs
8tVAEGNA4Lt91j5j5A1o33/3GvpBqHy4oQbv9IEXUiqcpjQPRzPN0gU+2rOrogd5OzOATcBtxV9V
Re7o5kVXGbWLoeCWT5eov6igWrLYw9BSToVGQgl7fqPJ8NlLVLjOD6K7nnPyMWo9peD0GuFh7Agr
L/czcByDVpWUauT1DsWre3UgEFbK+uJaismmp6WURe5ScmeA1JMXmn8Ako1RyAcy2ZcSsW2WB0/g
8PDkM2970rQKtgxOcDl3PNi+LMQPTgSsmJznyMFOsEZZ69cGfr16Ckaldd2amKd14c2x9a+2wMHU
Ul/6LOWThc+Ic48GVyZyipEjijv30vs7V203ptQ4RLHH5GYDneCe59gP3zXNwH245VRhTvDnziOQ
FQ5+18SW4GQltZc4UrwFgrYRrF/IxiLUTRsNqTre3Wsij9Egx7xPgkcM21/gKcbIL0oAW+4bNO+o
goG2ShblPReWVSG+mBFfi6xl9Zvvv31oke9q6zuoVZ8KuvrjO8B4KI/tZZlB6LOZX7tl2x1lUkQr
eeaI/klQM+W5Yo5tHaQgEeOQX1qPH46v1A8nNLAMfZgiZnrjAW0o6tATBJl1UcYs8AHQvht+ZMR+
8cw1oAxH/d7Cszo2c6hbsCB9aa5t6kM6sn1CJYHFr4CLrnIKHncFJY3YNPNtUF6XdrK0IU4Yk06S
0bnUGELsVDvnoOQrJSgr0PUewOgRANb9HS7pH0A+lMH/U0mc37f6YGlCRVgfUWtcQEX1Jd2SxOc2
MOz38VOoG+HfffFddyuXaiDF6xPQw3F8TyljPtfl2ohyn/XUYKDK85NCYyxAh1TY/MnCAxcw/ife
py2YKa4XMLstPJlqAxOcA0PhzcpN1BvGqZ65UN/rR1FGlyiucbrJEQn7rRFa7tcPT0kVF5MMnKss
R8O49Zz0T8cA+O78GhljGFeQpyML3O+DSAc52+8cfO2MFk6s4E0VJKka2ylyw+8/1vlHXfg9v4ss
iGzufWeQ/7218iqjoOHc3R9a2FgutUl/Fl/0QbtWi17ib9657Cvfq7YbfM3Yr0lcYPIKLEGtuhJ/
LXMPvH6H5gMzZnhdH9VBA9a92jHxe5W2Hl50ZiKmnzqdnx7khmSFt45IlCsUee2EUySo170XOjAO
lpmIiG4ska8FY7ly7vZ4fifmh6b84m1C6088dlkA5e3gJN0430pA8NJoL5HBPN7PIyewxBHu7qyr
TuoBX88AL9aul5LPmGZUQs2OuPRTrbOuXz0EaohJJ5vIqyRmWCjJqLIkpnTAILO83aLZhxWpmjV8
ojo5ngiIO3VVI10LnCjfbyS0D7BbpHmmSnMRD0LeP90HdlQUMul0wTxXhs4LRdACK8Vrmhnufxgb
5RKWheN26oCpJHWeiGAQilQzZLzO6ghMMsLyzZ9JY/OhRPcNpMjup1lEjMKrtoc08xqteD2sBk2m
le502+dlo1kKwGeaV6EOVUFuYaU7tR5ONE495fDhaJDfx+Hit2kz2W9xzCWJBA4JwMKfZeIslc8r
OGqRy33IDiqLlYYchwGI1BkSW70EY6rhtui03VwE1UTkO6QOI8Q7O/wdWFklI5Y54NMP3cw5wJha
HgvBJynPlNUo4vYh+/JVRLkq62buHr8zSj+rSPoIfjj5K7Y+gvZVUc1Lpcb1s6fH14RPG8MqS1g5
uHs6icqS2reTftDN4+1UjjvRjy7XrvISxZiuRzr+bQQ3ZlfwNT8ser7NbQ1y3hvcXfzZPsMs0JEe
/dogEBGJ76Mm5IWD2TfQDSVihHxRjc+m/z95Oao1rZzE/KamN6PtYkovHKQZCjRy4ktrzEbYWIR5
ImrY2yqfB3+lLEpC5i3kv51wFk91pn2CiS2u1BWMiCdu2kFj15u9cOZVnxCicXcN7C/QqTjbovXW
vXg6WBwAy0HX0ixGrsp4kv8rZUH6f3s7csM5uNNNXHAllBA9riON0AqsyBPpha3q2okxddHG8CMM
yVIgYXm8GUNZgSFPEvNHOmcWATdHli/0OU3oR7cdranoXIEVG1M7ohr0u+o5CnKa4C9mafkyiXIT
Fd9ifCHh/uhkl0BxwI8KA1OMUPgb+RhSNUhLDKMwaYBB+2hgaLtsgHfkb4qzxRU3a2pDz+rG6EW0
iHM6BHz9NIq3oxKg4zUtdgI5PoYUfEiFaXW2uG4b2nNZswp27igOm727yXk06kqX0mYEWOgMrkPm
SzYYPuh3WytX6Fu2qrqeldfJLaN5uONVcM3gNoKUKemJwuwQtVdA3cxl2y6aSnK3lLwj61ROPPbc
8s6MeZlSrWCGAJO1y026YtAEyQMYW+LoLsSJWFqG1nJP1U271uhaPtPZtshuziK/PYqGgU85i8Ec
S4D3Gl8DKJb64lev5q0QlAlv61O1K/JIfReyGa4UjiyipUW37NJUGSUXltLLrRLMHmQ4WKlYzciM
NaCIBphZqE08mD0KG9WWieAOtHFu4ODo79AKsXt1xFM1I2dAOmuFcOuSUO8OnZre1hD2mWW9CN4U
rQczLGvTA0VobEZjXRbGcp/qSiuBc4VyLy5yMhvoWGRsaDyykIokst01ryhWf2XZQ45g0XHtMLTa
3t+LowK5xyRkHzxXNpcdZCRbHTOkSOQmjjBvo2BR3lau22Q2FSTbRCrif6GxGM+Y5d1qZF2ORGIM
smq55dIm9oGpQAkjUVL/6Pn7yAIuJDBbGmJ8G0CEV/Q4HqVRvdOWQaVf5hAkOVlNczU/o17NbRzK
I3vvDp1sOfWYGDP6ngO/0I4LWEw3xK2zrdnCEovtM4iT8I4y1CujVJWA1LZRTh1Y33sFL5wnVdZF
iYSNGzMcnBjiY++RbYkMOB3KcZ97wowezls/BxWhCNVAzGgKhSxinlRgTUTK+Bp3QxwwPKf3q/MF
Wjm/uhFSyhBWzoM2Eou/GTxdj4Iu0gqHy+8fsJMc2TUP6DD1orbbO8BCMEYF38fgfMFEPUeTLE/N
TWUII2XrhIQXC62NikEK6/TMK+XVorws9aDXgVik0nLeZFz6IvaZFTloWgHBrZWSiDu0c19SrxxL
EjfKlcrU13Cxll3dQwRMnaTA7qtKQ/LJ5swWHGvLST7Q63Oh6zR7VYwaALld+16vbx0SIWMWUkpx
OHrG8iCO+WNhVd2ebUdxwgONiJg+Se7PjmCXyg8ETfn6gWidhkL/EO5UaP4N7tZWccjKGl/JB7zn
RYFtIZoZJWtrXPzcFT/SmNF9+qaTmPJMgagOFiqypr2AQhvqlAxZXuKCDHyGAqTgvO0Pz70z39pb
0KWawtxedNeHtfl11tm8O9+6qSs/umyeSi2lrwmWGck6Li1Gfwvm2+b3K6TlptJy+rumn9IgC0BL
4lPDnqkiB4ioUsiRMUs6zaCBQ21M9I496xDvtRixjCF6VBHIKI5MBl00i2JorUfzcgKIcZ/xtUx8
iPnMyGRtaiXW38O52LL54I+W/t19PArFL0pcphvKIKbNadnkeAlJ93W6BknxK8RCdp0/XfmWamFV
FZtndu5o6C73vzQL+oCDIShszmeeRIQvJ6saA7dK9oVPfPbh8X4v7PKQ02q9p+UiMbAxbkBhvUZu
Fjgh5Avbmabp0WaIno8x1oIJW2wZFiF92rK7f5J1QAw4UPZmAyo2gkwFcftIe21q8jQrOxMbmBlT
Z2AHraVm76mqKV89BXMj9mUugvTprmYibwG83AcaFPyaGSbmYEGpMwA1zORhQjAULOe4mUjpql47
xlvXIHlL1vYvJ+PEG+rGBauCwq9KA5+oeFUSnn06YVY9HD+nfMwf+dmJZoQ4DKVDUbIweFokHwns
2HJ2xAYbu/SdmcMy/gnYA6ZrpU9RdJZIdya1arN4OLYfb1DBBoqRW6JW1q9rkiBudjXfnCju4ZIC
vV85cGzLL14gcYh+Au8otE8hn/NfQZjcVVzY5W2RH6Mz5iDkDk/1r2YlHywXE4AyBgNi08r8hoZs
SXV7D/ABj0+oqtEQ4xjq1yJakmyD/DaEMwvqjc+F8N1f5Iubv52WeHLnPxw6/TGxP+/BW0v5ktyo
bZXzf6RaMF3GREyDWffB1dtNiX0kmROXa8Na3aQOYnQmyx1n/L6j9A/tfTh86ZRgXDqBieOTsER2
MV5WW6yqsAIPr28yIKE9nzO8pzfxgrqNkA3Bbm1FOggle9A987DXs8bEXz9H8E2JuDF86WvB78W7
eT/1rQ2hS2KF6lzKd/tULc/5Z1GaTvQjYMjEHpPmTx1MCVNL+A4f5dlM8tKq6+Zc5XVuVojwZLTq
VArCIuDe7ZosXVht05NSGXGPpVojFqvVVdtuTl9sslLeNJp7bREMvOHfR5ku4J2OHyr2iJyeLCeF
oIZ02DP2Re2/v5q9xPSQO5EmP1fOFZegclKP4/9vSCR+IP/X10hJBAkW081QZDDMBbtOiv+B1tet
5xQucsCSqZcOhNlUktcIT82gacJxN7yj1a6RTmJo03RGtjHzrOZALGQA5eqKwUQwmI9ABSelFZV6
MsjrLJ/WVwLK2tp03HLEdxMuFj0Lf7nbRq5R7k+aBjyExmKvbXVC37M+9LGEaOWycUK9rroK9jb2
awNIS1Bb5BZJPmC7uTcBTfsG5DkMRnPLNHH49tEggP3ChO1ZNxGtUnLLUBn/qVJIcz3HoMlvs73h
35rFOjS4Ij7e0XxWiatGY74nuAHQ0KHtDq+nXa9kEciiIpAn66JCEU2vR+OUREMkURKtlc+PKlg5
kWAsCVozyOw4Yd9SCHZy55ePXTRDFJUE6sULb9KI5Rcph/BqOeYNzQrnOPCw2vEiV0/De2VLOWTq
9CySq7tDKbfaEJJ8wfSeiUBO45CBvw2dgPG9/AYhD6JrjSDqOCSakQSx6Jay/V+EIGgnmo1LAhwP
SEaf6jxtdWFx6xu2hrIP75zn+CcpPgWykugXzd56Fm7jTtMqX5SHf6ROl3t8tzo2IT5qklTK36Ys
GfftuTbkMB2jLyZ6orvIQIlM123ocCatZN7GZMiCCML33pRhpmkHRj9BfwFUvSUubxoGFAEy4IpW
mKXYiXgZCqg/4i2sNc8SKsr2MQ5L957Th/8Und2ownUSklgXEXaZMgW4gGhsrZPR8obT8lZ6Fusf
shqqh19R2ZZloJ6JzKCQUeKHtg/1cQQ+7WMPSQrhQVu0mxfe/m/BI/vuKcNf3F1J1j2XGPm1E2b+
z9gBhW/LSE3rfgCpYSrAb08RsMzFUUYC4Mb4Ef3FMw8SuFHZgSE93+DuuL+vyT/KT4rSMM8yeZ1o
vLUJhKi2hSq++9j8mVKCQBzxTPDcrsrboneSGKwag4cDIvA4L4VGmJtk0KqjKYdV6yJVo6MEbG54
D3pDVxzB2Xi78RztC0i75dwsOo2i8dfWnzvsa+UJHEX8/gfL7e8cYOeNbzuRkNUTNbLvE5sW7jDJ
tzM/STrtDsenYB5UsaFfUChMTzu53EcU6vex24yBW3TEr93jgmo4mWFtbnFh+k4A//kAd67T2Zv7
k7ehkphbTy7VDaU2bVAiR1mvIiN7nVZcGzhLrsZiwc43LwJxmv1Y0jx598sJ4pJLZwXWjIc1GXol
q93l7kNY1QyT6D0gU8XVd8B+qbjAqNd7R+eX4tcxeTipo8HU+jjm+UxSsURQItkD/Pgw+RA3q0rE
og+KS1iQAnOpk4RDy+MpsNlQuMI9Rxx30ZQRSE3cL6kRPzqJzMnKR8cue72cIq6HbDsqIQb4HKKZ
i4QuZFOEcBsKlAe/Oranoygm+BOsOHzypAtfajhqZFQsmHzg60D3BHbkoyz6OWu97TJuRcK6adRA
Tkblo44PuvOW9olxCt7Szv31CLUG3nWWmX0L/pneKlg14e8hmhgn4Cnw7mCKZCV2YS9PpD2hwoYb
AWAjDS6XMzBgJvDg2YnJ7BcPu2jjro9DGER7tpsBs1xZE+ZVtARish8o+tG9X3GR7i5NNa/MveVq
tBfa3CsvZp39Ozf8fhF50IuSYWpBxUdnyI+8lr3uX+SKwWEp4HlJVG2retHqZWNA3A7fC8qL+mea
sgxQIcHNcMeqYEGL6arv2BWCCaznTDIiBoInP5DvrqsalrxUSkVk/gEhaTPdN7af9UOVQvuXgYve
8AWQVv5jDOVKw5W45ANnoVyN77LldXZkMWPArU6oAEjWWj+u+B3mvmKrXfLYZTiGXcONONo5u7uO
4k3RdDUYFGTzhkdK/IXcnthAmTnMtz5cNqS692Hr8/ZP8aliRFrr1z1M8/nXpzkt5icR1jFHoJQK
3cvEUE0+ILWZpHJ9dKyQVpETXKcfDE5Knd+N5Q2VuFgkpjFwtihDkOGzUgEDseWEPQHtemOPXMAg
TpKNg8gYGsGpJBcNr4I0fCdX4yahAmg+JUaJMuwlODOau/NkNPn4e8CoB8YbOUHI4QiWX41WeNpb
9AlQGYAEgQlbBre6+gLYrJEkKpUleSN5Y9eLAifgK+Fky205qzi5ut637/u55uuz7/t6RKw1d1yx
XGOk195+C36MabmhHbPHsEIB/g9Gueixokpx/GzwsAimEoAS2zBUIlrAWOK8AFmjLKp6MH08wyxp
PPmc1aglEH+Gs8VS/wASqKQXA55ARbLpDKGbkX5K17CGY6PJopCUX7L0J9QCcBC0b4RrJxs2e/jX
SsZon3hpGz3Kj6ii5nCUhm9wCXfe2fHJtng3jOv8Jr/WsM/0GnDnL5rrq8o/ON/HwpJs6neH1CVz
RFcMOH1dJDLV128a5nkH2WHeOc7K/2WAFJXrPx41k2uhQ4ZToUqA+2QpNWvWJld5q7cTGlf1CDB2
yHKEhMdsdIxIoQb21ZX9riKlVoJHj9nndye4DENuBA5fh9j72uPtFlvnRzdOo8rN5G7pjtHX4QsU
1Qnym7B0OdHRU03ta9l/QUFbKS8XC3Ugd1DmVcik36NTdEvhpjSwMa18nAfbtToENxWMAs1oHaZN
lKZVW7D65t+LxW2e+PiNmhjNerBM2ToMYkKl4g3bBYVuY8X/I0GWESTgMpWb9lL6o5QTvwafdCD9
rXrqkzlpctJOwnYmAi9EGAhOxZmG9HPwAYTFCiVHe9Vkr3mZSHWM/sfz4UGdTngy/uoJMPrm7xC6
k0rtZfhJ5mjhNRSjrN87XzrsiweP9KM2+NzJwWwBy5X52WyfMni1y2/bC2crfxqLws/yMUrwkLVj
X1nhSHNZAqi7yPnV8Fjj1JSX67uW3F28mC4jlMvay73a4xYhaMK9MrrR6HVP7njNve1ACgGuqByK
j7bQuWnbJkBgN2bFZTHoRwFRRXx9Zs6CeV+2Cisev3VDVhJoe00Qp5gwjY0AJYT2mShAAf3a9lJE
tDAfPCX/l06R5/MDAqvF3Jcm+QbXAiPjx9NxPkKCUEVKXR1XsYbjYllkcIJQr35wMGLxLZ1DUsNR
yqg5sY8/8hZPFtLJnRLRQKpay9knKmQ7ctwL3kt0FPLicipHJenAN7hX0El5aKCOQSI94T0lkx8d
C8yH4jZKRB3x40D/U35LcNkAoQ6MAyBuMmO75Jo3V/ZCGyRo2aCEGoF3QUaxKjiIfcQ9zRjq11lm
v9pj8TwSBaC6Ek7jY6Zo8SvSaLbOVnxX84s97GDUX55Q1Z2nTOgSRpH6g/P0APPMvMy/BjXm9qKP
i3duo9vE/VPEww2F9GbuK57cLm0QsrFSsPirviR8lwkPOPUZBvEr94jxsjrxQ0yKeKebWLXQLM9E
0/IWGiMmEY6iq/v35lHBtYA1XVyqgZv/tEPPi28g3IvIa75kAYP5iWU7dMdBNs8CcsSZozeNGqGr
4FY9FX7HP9EokBnJmHI6+E/7lRG27+U+ZqdB7yiCXYvXBwqKyUJ3lT6UyQs0GyyQWTExK0jUnCrv
jImgIIgJnXdKWsonLgBy9IBrrjtcUo6K3kVTzz4JzFio2HKko73ypH47xZx3GQ6fyeYQOwUgxSv5
RBF20LCFdo74c4FEgSWsAv9oXl5setgwAdyONdAqqc9hQUKuCuuu5h5fKHGEpwTiwI/Y9L7QkXTV
sq5y04lDDvIzOeDyFDnTXRmEw1dM1gratmXYDt+OsgY/mkLwQI0zyrEql5iptY5n/qfCVzpi7hIf
/34fTs5bJS7n8IaIEEsN8ex61OXayyVWddTokKMNC7iaSc+rW90fNAyEAXRbHx0zhncOxVHooSts
H4mcvFujkRmCoKUrhsYJ+1KKaVk28IcSfZ4mwCMFUNFarxvDTQBCws0G/+zD1N4qdCyLUtFhSzBC
lvuqy/q3OOoUdrkD4z0MMNjfM4QzlEYdQIuxJ3/rBk6NbVxUX0Wr5qVJFR8wjwUAEDDfZ5DRbnuY
gcxM4wvFCsY0GUytQHNj3e9LsPN1OrmDCjh54bX0I8cM5HisHwKrB8UjSjjdRboToU0yQuaXisBO
YqpuZTS0FdQD9GGcF+wyraWt6i7V+CwSOG+OymI6izKsPHLHQ5uknNl+rSwuapoDg1m/AtjVou2W
D6oeh+8G9Ybmrhn4rAvvk+iVyHtl+rj3pqL3j2vhLc+d9rkJG2kOfWXJRzh93/vKjQ+iDu2wxwEn
56KSMQbeG4dz45K/wE9wclgoGBjdYUNTXlBS8BdwbSfDEN7uR7Dp4BRUB4yp5ddlscs8Rrqywj06
ALUhir+k35yPg3qPJn0NgvCd3q9UpvXCQrlnA1oeMrBWmO/wcxGFcasggEub3ZDUvR6vYNalPFhe
kVUYOWkQiITmt7mr+3Ww0FmLoRQhkgpFtAChC9ETVqw41mzg65S8fcpXw5WX/j8sXhCnpCHhHawg
oEp3pmzBDM18FsfS6YUeWX/6KwWE0+bY9L2blFPmiJ+wQyEEjq/qM/jGTu4mHEljEyePht+tlkKx
UQ7XInUIK7B4HilqTl4nOP/jBL4cj2lv2sojBDh2NTsGCC+g9OGsSTBPZxkPqGSbEJFHA9RfvYG3
Ac50YcLV+kg/r00+ReXvEWq+luOkzc5rAg3vA9zvqTAodTj5LPGWku8WWs3NXEcWMy4IC6mcTAT1
s7Khhv8wPU2gHGJSh7ldQoB/pj56S1NH5P4Rs/mUvWvK7P0RuYQ9+SmPmG8sD9MN1VAomKbncCw9
ISkZQs4ieJVu1vZgIFuAiTe9DE+QjXjg1FO6jtJSmoyy/92g7qxbvRUdvM53XJlDmY5zQ7Rn2YLA
8ubXd3M5inJlkM7AxwNDuscLcSVL8BctXN8sS1eGlaF2YwVOwXcV5AP0cT3O06Av5DoywIQyzDPF
PviXhQmFzgJSByb5PC1gO9xNrhBQCmlK5GSEH1GHktz1rOXavsdqkYgUAi92JkiJwdLyrAOElu4c
yd+i3ZXaWI6mwpUPrnemEqQ2s61I4t354wSMtKFOkB36Bb7C7/aJa1gR84dw3eA7ujMbUaWq8884
D5KcOt0LfwX0cCts4bwVRdqgs/Tf21aeuCyWk1sVJbfxEkEw+GfKy5df+RFiIdqYST66dPxeQK3m
xsopAqdZKSlaHX4mmSB9eoJg7IXnZiDS+MdxHSWcgfw5DmdJIbVFXqmRYs6/O8cRf/XQX779eayM
GenSF0EiUt33SzkpmlI1h8pwq1mePdX98EWK3IWar9FR1D7lzD9yyUhdMoDVRjoK1koKLK/Nxi3o
QwbjFR5v/Yi5vtbzM4JOFFQzK8NnQPiiuWH73UP2gx4dBhI/boc+z1euxBNvn08adGdTRUOY02x7
4IXrFZqMezbOD9mAHkDylPsY5jJV68ThMJJ34aubWySpJ7fBTOVg1sz1Qsc9YqumfgGMsVfLd2TW
ECKYt2nZLcIxOU0ArHRlgGJ01r2R/9MFZP/oy9/hXHXt5D/XWuVbKVo2NZeRcqYTiG8rkqe1goVj
KwZ4eLZSWJTGI3bv5ZuOSAuDSJDNPeb7rknekd9lX8ybJ5smAnpC3Av/EhPYbf2Me+pI1d/TDYP2
WCctwKmHqwaHhZ1u0yt3s0hW49wleV7gapz+XpwxNQIi6ZTGj/5n0HesOQmTrYXoXuc+BjN0+8h9
MOuOQ6k0fDs62Gnz1C9gBtniUd93m8Sb+h6ucztO+vr/NVVVh4zTisA4ZsMwwZdNcCNzquLvRPUc
CKDWrJ7BgeISQarTF0kkFQfl07SqEjFbgNQD2r4Wm6yt2uBbOqDyf4Qa/zTqcxLR75sWPPEul78/
ax4Y9+rscjCTpU/n1VHM9EzPdVnnKEWw3ygaFEf0CuoUROKB5YkymOHxmOgjuHjoDBRKvBi9RjE0
HPuRxKwgE8kKQHsq475YlRzD6vVxgcHfkWwvKJn35VMnS4x3x1J9fmvgWPUV/r+Y5OfnkZk5EAd/
fMM9K7WPN4sDX454riVqEM0facoKSYsbgnicR5x0kgtqb+PugvmuJZyebE91TaiJDESuK6zsKr9I
Prz2l9KHX41KH1yWYmR7ryvWLUK1s9idgtQeWevp0Vw9wnl8ifNP+yQLYIpv4ifh7twN9LfGFulC
SkqPNB+cdpfQwvYTqZn/OsVonFqrY+beNX9zNPyWZ/1VtZpJRT8XbPwGIinEldXQdRxeEs0OBGqp
jcj6q6IkgSl58NOvQ2mCnjRNlJZR8h3+xek3d4Z6N1HziLlnd2ItbpxX0x+n/1iUhgyelldqhZZ3
TPO0WisXuCW0hC5/vckuA6ynmdmOG0c3rH44BcYfsAY3hcs3SUSY+/XJS09Rm0VFsyLJVFE3wUcy
Toj/MPwR8Me65gyxwNTbuhzNi/tpLY9cQhLcKOuSiy97NnVJasvJfhhHu8ewD6P2vQSZT7hi9jpl
uqBXGsc3UPQkNG0uaXR5OO3+JscfPGyr9q0T17KSOA1tbxWZgc/fPVOmZyWgXP/3sU/ELq4Bkc9b
V90ME5hWumpIxK+Uiv5oolNOPUUFtDtLU1dTNUkbq2AOi1pYXRW0qKcr0Fsj5YRcKQb7/Wzkkf+k
kGWROpRZz72BZSKZyMIxYJA+01+rdfSs5f/g+vB97hYaNdrX907nzz6La3WHCFYhHlyxP7Gn6CAQ
qTsR9SUNYhqVOa4vEkNCLAUaL/6A7G1SaJPRiCMPuk35f7l7h1hZX6okXnwq2+3vy8zns43LNL2q
I2hGQd3tr2d71r2sFWdDIF9IkLsInaXkRQg+6VRHM/tqlIbG+r22mxdL2kz8wwFqOPnePTe0p45i
rxhsk3edYr/pndD1Dd0ME7WZnY+4PFXbB0ZDJfBqvfDAOdCrpKIK9YswO4SAQOmyHgJDlq/q9j12
n5sxlcEGC1uFC2LIGn4HcbqVonD8EmwWNMxWDdYUPLXv9CnRBFahCBFBSpgybF+CI9AwNsEs05nD
OWQFYL6ZUJ1W4Y0YvUip/gX3JY7m5chmg6dy5P/iIoVk3btQKsbcEfhgn9k1mTyGz0K9X1aX1znw
CUFFq/mxdvdx3nA5QWJNGmcP1CO2Dey3ZSaXbpVM5hqeIqjYPSsuprHHtU31IL7OV9Y++U78Zx4n
8TyRsn5DPscEvQRN9lWy1W8VxbnUzoNDXIHii1kh3gfN569PLNZ+FzC51xh9tKm+IkwAGpqNBib/
yckBY7S4+VsW9aXoxENGo5xjBPA8+rKy6vvPhu9eFo2A2wLk/4VaEmFfG/x/zREJJxLdNH3S8Dnd
dRFTMxqOJhkVCuAFBz8GgprSwRV/SX/XDIbGS1mHFHXOC5pCAmRW2/xv6LM1EDPZIbrNyn53q31S
n84/lTFs22syHCUNETxIOiXrGVPL4y80lkV1yD0JF7k85nnSEapQ7f5/mCtgFM5q/IJibsS0nVfo
QAD99Wmqw6GBhwEh2gFi10mdDNe9LzJqEQ/UQEZu2qOArLSBWnxHeRZGC1/1BwxsKAeZI4g8bNRS
KzrvvpWOviJcM3/t0YnDFNFLGSBsFQOEm9X9caYifTK+Kzovo28r0+ZWnH4GYwE3PZMil8uO+LIh
Ir1Tfk/L6nA+ypRPCMB8G0e86wVkyd+fVXhve/as7iUg2PEYr9mCy62P5EScx8RhT+3gZv+aSQX6
RFhAcgrKLdiniZGLXEEUV4xEuNjQL3xqyPcoVbYzM72If22s89PR13Ozt2MA9Gabwmx6AAAeyvM8
EOhB/HDT6F2FO87RW5OvMwi1zwpcSKBOFNW53I9e1YzMuNFJpK2IYGr4oEdDGawxTc8J2j51zNB3
EmmscTYrz+9NfMHLeJuZnRfjJTCYE7XaYzDfofVy8nvaJ+Z13/sQJYWNWbQ9Tmnh6h6TnmlSCF++
shZherk6ocuX73zbZio4Z5bZr1edHPlvN8VTvIx8clIB6OtXxowz1qnoCn4WE/X49jiepgu5+2j+
2a97/ZNKwZTAxxfxIxRolY/CfUjaLNLhcHBADyYjfhEfb6v2y3ekZs5gyo8jRzSPxv9B/1aUrycs
hqVX5LZwOf2oDe8Ko3oPlAZsjBxtCAZGZ4PPaed6A5gP1h2KX5ozpFmiyfYktcVOOH8kohztAPkn
Hbvcv0re9Y4nWiGG5dyQaD7+8YHqKKb5QfNg/BYKqEO8VGByWX1davc6dN8NNmbAQ7tFFBNQFbFT
yHefslirSN5d1olMChDdNJttByTJOKJCxVv/grOswk4uDVvNT2cNQLnVpw7B3b4+X3tGf8Zku8a0
Q1SZFPyOANIh+FzDmBw2Hpi2jaOk430AaNSGeGdurx+Zii3JezvwBHhDaGaauacd5btBYAzjBKyc
b4clYdgfWsbPW9xi0OxF9w7/rIJQvn8ruUlcgsYI6KUTUCONUjPDI+GLVChha0BiRlm0UoHMJ64c
Lrxcpp3DrhfGzsV87Xk8YpFJVj1cAH6WQQQJ1LOjWr/wZc8sVE95DP3w3X52BeNka7gPaguyWB8r
kn4wXIVPJXjB+FvbDMiU4VbJZZMxwaqW6SaKbSsHRQ9vUEtpzieMPdLTW47QI7rf92nPVwMKvukZ
6NfAfQAZLHVM9Dd6V21QSghyMddwKPzyXwKdZFSN11vi3bqpBWWgR/y1sefwdlIRv3PK6tO/epac
k2sAOWJnT/70rsZU6R1Su2O1F+WSO3oVaSbmraW4MlYRrx0YD8DAuxKqmITVVBXBPTrRdepE+eLK
Q4ckf73yt5Nn/ZQkWzSgaWBFac0jjZ1WESUlWBok3y4Ymh+M8b3bDjy5MC4IlTWz6BgpwYr7y3Yx
5OSajPGtXmpanf0XZ9HPIWygYTBQ3b7vzJKZoo5gNPgkpHWVuS6z6kNL05408YJGfSrY40bSYsjU
w48wptkyM3PXfPIplCdZPHHVrOPKFyvWQqsuNx2TtmsUFguco77B3WJ0bmQWL1Ljmkl1wVutGjB5
G2jAcjG5YtXsVC6z/YPpHYJY9WmP7AfdvR0yl2qYvPCn8M4BFIvDczOcEGnyO58jIif6EOXzMZ0U
HRFH8f5U3WvvFRP4BCELeOcrdww+s54n775TX+3NguUTe3ZrDcvcXXdslmbfyfMpJvw3rDBOCavC
CB1A24PLDNKdRfAHgiwcTYljDoiTB0jeNezTU+s8tbts8qgFxnzyb5v4T14bmjN8DaxSzEFvZ6y0
hRlJIWNUknf8i2CegW9HUuzPN0e44CJKkSh6VqBFgtrhk3thE3m6+kP8itUQevt/jSy23tkbIVRo
47U31Cd3Pq97JXOTrYwEcyF3hierJX64nOEBOhh0xpfrseTMm6+Wr2d3XLnfrTvL7F+xv+OskDIW
2Qo0oRMzFV84hXxXRvlxRllCBZB/wKsSaNrB1wvq79eWJBo1uFEbMVc35fx3jTtCrkRIBgJA4b3L
Y/EVHHGHbiDNvS3uoDWUSqfzhcNog0PvV7bR5MbJrQbwHXTZWlSJqDBXlSPcCXbXkUo7mQROb7Kb
Goymk3wi8kXWTSL4nFcSNGFgmlGW9PM5bGL/suzXuZBj5Zoo1d0ATYPsaPtBdlWZVMA73rxEA25C
zU96X81IURwoh+X26MH9gJqSiWSDH3o0OvZ4tm9DwXO2d57fTZjSh6WPlHCtEHd53WqCR3QyYtYx
zH0uIY+zlRZkh99CUd2c/xI1/phokB+mYuTSjHJzCphn1wONIBVftIoqTyGEQxShkuNpFLUYPrSx
Dn11ose3Y9CqiuYECjV7IqMmiALVmpvyOxtmhtn+mVV2utPUJCCOoUR5zqYoJ5qof+Q+pBGOb+CG
7ZAK429RatTJPyIlJiVDgiTNQNWyoHRPj37RO35X3Zn/LWz96yTqr2O/k34qxdkykjh85P9IjAtU
izr1raSUiYjO0kbsjfr/37uKxYSgcrRdfC2fdIh0T4w+u/9BvxSGAS8ahZftoTuQp1Q67VlSAEvA
TVh1ywu1/kSsCI8X0L2eyUSg9SBnMW38YLvFPTdWHlc3r1h8mLYSGwzp6AVIIn29MqlwGbQAv7vY
EYOfet+UeVHpYBBa3aNYIAUcu+A8fBab85mYAAXozSXsT8TwYw637nUWNFA8Lu7/ckdbNOKEObfU
deOf+lri2q+bLmsvK2d9Hwh/w0yItHejnsIoqHOz8qec4O5aKFPIKc4oUQ57cSE5xp02PxQda+Iq
UemIcpFP6jNQRFgAPGgmKmPGhBS/x2WSxZwDYj22Nzzu4mMGTrbWh9I5BZOLvnSY1anM3D7T9q2w
kePaJgH9jSFClv4X/jnJl+R2i3H8TJD7aOzE8XgRviPH3PPSeL6IGl+dKwUkmcyJ6pUhH04icDgs
wt+A5B0DazSffkkKdhFZsbgFk6y0Jhear97jJfuRXyk2o9apH4SztMnWphOPNnzQ6SRkA1kU7cW/
ldoSv6TEVzG4ghH2CZ9JS+autq50MGUGdTR1r91O0ljGd/Xs1DiJzvWt76DguNxN7YXHPbC4Oe6H
xLPvDACvBgINXiWgG5BVyqDvAtzlKwDr3DYGZ/I02M3m5M6iBTmCDl6mFYqpLmb8RbDDCqA1TY4i
DSvOczQtNnsGc8/SMkpG7TNw4HxsCwe+FOOGUnUnLRRUMswTXIQNppA+Ot3o7HkR6ehPV4OoyQHh
dvZMZFJG429GNp6KvyjHfrgfLczNEgHSfc67omITjo6pBkD05zlGC9d3z4c0jeoRukK57PBCm8A7
tkhvGjOA3f54m58Gb7EtYf/PbzSGb70kGEwLEo9DfKh9DrDv9YMM6/4PaGBgqApkOCvx+MKvAWGe
BbVDpHF26sSrRohMWinLp43G28DoKMsUnqluKFrmy3tyuCvyc5rN4Ws3K8TRc7WkqNwpW7vengoN
Xzeaz5TPKeNCW6cbpXEtCk4sp0QMz2Ql52xSQylF2JIlPZHSZzGJ67ythasapmYjbjFYyD8t7+3z
ApP3HjA6ytQMDxP7CA+oXwBfsn6duqJGHQQClBSjSLergod1snOSrrNARdHlWEmsoxRawEOVYBrQ
l2Y+0+vlRUcvzMb8cQ+PxN0mji9FZAqK33xPBe9P829janme1IdIG67LsBh7mqVcDVNq7iAEAXN/
ld6QlIjaK0GNegdtBytIVk+GKSNO8JRDZH8EG4uLYzA8DV8g9e4M17tETrrsUm7WHBkRBu3at+N4
ohkfdKeah/ixMIVhovkMQL8J36D39nPsaneokmSPYhpyaTCcak7CB5FQuYTRGQ+Gg1CukaOUjvF9
dPprVeEkUOuqBkxjyFZl8qv4A8ICWbOs9CfkFhDdE95wrlUMdmTGbAsAK4jLz/2UBhwULwjVHpxS
VyycnYw/6rXf45fQj8RuYiBkrQzs2N8qu0CFZdTmmog57FGXM99UQ09nyoeJ6RKfN9qFZbyneVRZ
L3WaYhWj1gqBiHehd7zP0791wLWjfOKomsS3C1pGUuo4vVYtTrsa96/x2RMcJrhPVpR3mfTvcjkn
MMDBigSeuXNc2/qHCubO07GFMno6ZGlHtnJLV8bIX9GqphINR3ouMvPYCh9aIPKOYjolJFslipuU
6kTd/Q6h0mtGKG9VzkeinBE/qtBV7xlRFG00Rg9wmGHAkxeqyw3yKN/70w1bEWa0MA8cMtqdi1bA
LFBOc8f6JsQPGzqxf/M6O8cnGOf8fObU6L3xsHw6xU0lIlpxLZbluNfucUSpQWgKkH3qqHUk4gdE
EzSHHlT8wao5JgcqqPXvTB8cwv3G6px64ntftgMys/i9IyQzFZm5c6p/70FeULrfd7S9q5hWFN45
8htaAoOHty+knGYXJjwvnf/rVDjH5dVCWpHFUmkzpo4UR039NgE6XNGpwQ2yrfpj+kW1u4+zpm3h
mcn4jfNr9uOUyIOPEm/sHVKMPqeNqp5k16s9dShPeR+o4Zvj/ZOHnHi5PWnjKxl7gnwpDMIkrFq5
lZNHzVOohjTHyARRNMRXFlEmlJ+l0mMvKLayM4VwA9FEofSHvLKYvNXbQ8unQ8U2ufJaj/TBADZ9
EyAI//EGvu1FwRPEW5gHk+OqQVESx1OpySKzB27TsoW9Z3XxU33qK0USKCQOBsRjZ/lq75Ujyyk+
I1Hp6YKjESJkT/FCeu2KWDomb+76wngLvdGspx98Da7qZhBxVdOJeoxlt+LIj6C92fByJ9a6nL4W
OiYO3fU+CGhlttwRPDdCDaE+BTlxWFm4WMyMd5l135XuAZI9Ot1c9/405puj7xXutyYfb6g3ZUto
lNfx2jd1HiMHD3tImY8adplTiLc/Visg8QGbN5rzJA+cceSPsiqcDLiZbHmzvAtergGMuBzJJOxP
kyDIi/rD+0S1n4LbTOz8dyA9dmtsupNmn3AydrLFlmrCJwq5Ifb9efM6HcCmT4E0nxt/14UayPAP
TnA4Pr9C+7wsFprUBTtkI58JCWrocqFCTeWBEb7fVeHfnjXZi32tIrkxltIWtmYV42/7ijEdsCnd
woffyirnezFXP3WJekOmI+UWpY25DafGVO4O3STDEr9WF0IRe7rPh8IojsGahe9LPQTUXFPZqq0y
Yq+jiTgO3538Qiuz+kJjSefn7GX4jopBRs2XoGd2ydZTMMX9+2Lg5lEh/jVsgLuxvRXaBeYcKWpf
2lSlEZSrjVneJa6RiZpofIvi5zJZ6mBgGKtQkfMpRCH1HK4UGSL36mydseDp5saVC8jl3I/FoqG2
qlOiZ4mFzeCS4Y+m/pKARWDU7kz0MX53qYjVL+UUhoSJnoOSiCPGfwRQkR2qhzjsF6oBt5geQokG
gJn9inNCUBsz0F4XYwUT5VYI0nefxPs2gOSJTlZbMgQaRZFvnZCpNllsUn+hsb2O65kKJCf1NVJz
wC0ml7MbZigtyMy0lupI8qmzz0iEQ7ATmTm5BPjPkWgz2kIeZovjz+1xNeb9C2uuu3j79UilRobr
ISN9GaLyt0H6JQy6BMe21bgVmaBQ2bVppMR9r6iKEryMP0OvvN6N8JpM5R9zYhvC7tyBlUMr1hY4
9Ki0OI9ZVwqfAN3i17jCaQe1ZBKVOZ2UGViQz8Yu58+nNpoA3hY+qOUhIxYeagWIR1fqmBp87e1U
p7jsQha5h3gvRsvFEp2ywz/Pbfu9vA2HwNA3xIM5FzqJgxOLyoJzsRPPVgH74FsbMNwvt4lC4Xne
b8PXBOawvzUXBbFcd8C6tP5I6iPswoKf94MfVgtc0r/+6/V/YFUCtG7USwxRjmhaMM/G+tcq27Xj
EhBb7zUyv+BuxQmxja0vN462YLR8n2BtSVRDLr+6HFdO0uIz1zSo/tShoThI2uyF/tTzxkGi4MSC
tjYMH8v1SdHAQZY8VW4RWD+DH8vbTM12WpYjR8mA1QsvY4oRoc+RG8TZYkJZrimJmEWSWvKl+z3h
Ccwx6jBR428Kf5V7G8pQ+g+UNiOd2TyR3Wz6KjOqSvtRGU06V+e/qaGinSC22hKI0Ee0R9CBSX7h
1qr90S6wseodM7IFzNiHnsv7h5vANvhhDqvpLlWsq/dA31CgDYlzouz8wgh12aGZzl778lZX9528
JtgcyZRnO3y1DUCe1x9r0id8e+PdNWwhd/Zr+0BozmWulMr9oSkhVNICD7STz36MU4qFtEjg4zJj
6i7bCsIl93xtJdB/Ml9FlUPGBsdqpaWrhHjzvMeKzPDbIJTqqCl/xjWIG4KkRIzK68K2l7yVXsWp
DwjyejaodKszjGON2ilCOPA3DEV+jYi3+7albKF09kdJyVxmyd/ZxaMqzUpcyQnWMTFERx4DZrb/
zebGnDWL7d/ET8VxyPsurLgCawDbPuposxCuJ4O5KBgb7X62V7DLjHROVncd20sQ+JO8wUZTQbvq
pXFWUTxaq7G6b1KvF3BSo4oSf5oqiUTzuvC5ICnLHm5QjCoF/EugqsqHAUnvj+FLgNKcziZFznwD
IYt4HWnUW8rY9URGq2imrS9r8auHd6Cbz2r4rcyzrkKMiPefB/m/zlUSBmtq6YyEjIxSqvMjEx9l
srxYVIebJn2wpNw3gW1+gbhfbMWIfpEXLPB6lYmvuVhujBPm4QV7dreiwR6LcfRsZFfeDPmvv4Ju
QCpUzu1T6oUrDidvTXXfU5pY89ZcUz97RHO9nYu39on7HexSSxunSrCPaAZuK8jvGKvzXO28LQxM
Y780B4ttngh8U2/I9noViMwgQLVV5Z8Vgta4cP4LxF6azjQbCjWZFUmAY81EGrHRZGIj3jTue6mN
3zGiim+uc+2WSZhdAOymZ6O+PFGadGylv/pk68uzumAf9MKPpXyy4JUFTJf3Ex6mYxafAizhD/zv
eQTfonV3Y1ZVjHRSrU3muihZjllwyzWuOQkaixMQLWW4v1uZji9FbhYYDwcjwhf403iSIBxgAmqr
/M27q4mOVQ00oFe1M7nLfU2+LlPUHLYb/AiBdgLuOe7fJN56M4cjKPragRZtMppriXj6jXPDA8b4
urlTVb7UNnzKje0dTbvCnY0EcP2DfZX0AjJNXwQdwgZW72rfs3ETyd00Sm5iOGhs3YBXiFp4cIxi
Cfw2+9B4UrUtaAk80h5CDinMi9ccCZgHlhFWLISUNoY63k8ietHsS1ef32naHQGu3ZDtG1vnzGuV
tRn3GubEBzPtuT0be0NWghdL4vmh5rTPYNBQxnib6/Oes4yzLzTFFaGCRzxL7rOoHZLxCQfzxfE3
c9NLN0x3wWbBQ+1lm+H0LvPNz2DXQ6a4chFy8kBzIK6d3LQNBZp8CJu9WnK+HhvvL+GFEKGfEydb
GwNAI/xe0NWKMuT+bSEoNDFqhmYXuxMZp4Cm7OnIDd/itmuUCLd/AEGN48ZzoN+A2OJGXYupuP4O
HgGYztDkiyYYQa1xxhaDMR9lv/MTrpHidF4VyibmtoUG8MNorEEm+PzkkbzkciI5LhkE8roPOWcV
CuZKicIs38rIGo9p0gBe9ByGTZIdLV0OKr8iNb2r80fUblPH7mOt79EUGfW/uCGxAswmmeCMWFFU
apis/gu+Li7ISfDmmgGazf+TN3mUVErk0UZC0LUm/zaFsoOfrFRFlbB1jdOFSHy6GmPYheO+vJWv
aoi72f1O1vd4Zf6ztNW2BqC1McOEQ6rUS4t14LAanCqrcatkWnN4s/om3f1X1VjH1zPwYVO1Jbhp
lKlumGI06BqoUszHZGzbjhhU4o/c+GwtByoJrPFCJSE1Gzb1KJbHT9E5GpKV6KJvx4lLQUtUWD0C
vXyvcLIE78BHpOrTUmC+0n0N/c64j1m/60thlwD7ec/i+EiB1pvnXBWKv8qdi3zDl4/ascAgeTBG
QmjJrTuTgilJdS4b8QiZ98QI1HfaBV/sislnGke0V4UJSoc5YlCv8th/7OMjcLmNLcjJvUB+5bvg
E00OgPYFkbaXwYjMqqRr8YgQZ1IC0aRHodJW6oje7bPgzG+v+JoFvMa0fLb4uZ+Mf2tZ4C37EW4N
MnnCpGMmUqrrASDoZwGPup3+JLru9oQXpeAjyDLus1qnRcRdHKQyYJ9HQXM+v+81XVSCTlNdMRrm
bA3L1aVIMh1/yqGKpi46eJRgdN0scYxvDO8kjYJ2Ohh5Xu5zq6ESXH/Qy3O7ikNYQ7oumnkY8I5N
2yMgoldpFxV+PqxUtfHg3tXVVC4Y1OI6yrU8dzrJWK/Kdyp6mmkTbG/I+RDzSjQHdnlVYCAnQmEj
095OjAza5k+KqMQDr4/IfXw3mBmVkocR9U6VPG0bONTreBPgdBp1T91l8q0hDLjn9fdj2SjF9/oa
c3yEd+BFXGYEqfMAuXJkBlQP7aCSFBDaVgJBu7N/ne0QtEPSFhpEm7DPepSsHNjthpWK2ciISwHG
F6fPRL4VpTnctyXTqot9TfglMICeVrw13SUGPqxSuZdewWE6WglrMK9i0u175QiOURwBErmld05a
5+8fNakigE+XW8PCOfbt83Baq5MJTLa2+5FlD0Cn604g/Wie0tpXqmckYI4X4Q1tJJYzeKiV6zC4
NBGQ5oO+xQKxttRmERUc0Z7YEfL4pO+/ghlTP7RzmK7tRz7cV5bDE4k0XguO3UvJk36VoUEGjoM6
hVRPwtmDVCJdyPyCUeuiMjbS2Lugzc8GEeb08Uf2fRwTw94+Tal69uCCPV173CXzY7Uw8VvIpQaj
mGS9HoW/wvGDisEcQHlG5fD1+oow7Sd5+jyDPUVSCYn0fEQcjTYfPl9z64WvXkXEhdcuAsH9zewp
ePlWh6Lg2MSLfKFSGNzhfFm446aCGiNwJPGbE/geWzb3H4P8mhTLd2iMXGMehKpPB9Kzfh8ta/+6
qzcW9mHfk74lcWWhfhMoLeClwLXSVJtKuiH205SVmd863jmyiVq3eAGT8zgXUwq6G4Dtor3r7uhG
YVorsr5XE0+0MaCXZ1EXXnjNVXNpzSYCQ5SReq7pFoWlKQv492P50zQMk0DNKggwfZBEKggzPEtJ
gK/SVBkiw1503KYjKCL/5PBDH9/M5zyHw56GvQCr0oMlHdropySJOLaTlSiOUWWJloKWQeWfDS+w
j7YQZrme6SXcipR4dJcGtU2r4OmBz+tlINdqJLlXw/7y+3g714kXjtlmfl0Exjvietk6ZfIMhCdP
/CBUOYnjJrqirLzr6nF2dxgTfgqYlWCC7naiUCJXKTFc42kpc4+Dzy/8c5FYnF4hWZl9d1GQZEWI
nC2MBXLm47NddiGok+E4BGHH3YQtu386TLQYCeRqI53mXsXQkHiZs8dIQmM3OwCH87RWlTxrt2Je
gWRMZwrD0wSZh8d77ExLhTwYDDuH7EniB1i1JsfbLehSLA4k/fSTmPyWfR6hVH2z/0itG3Gc0E0s
xzwMRm0loT0KeqkEYAcDyxSF0tXteETMNqZ1Wq5qGInLh/6nOGfmOOrDo5bZNcZT5H8tW7zCo+cK
jsR3pTCx7pZt0FJcwGXhzoVb2xUWcsUqjzZq8tMCYIDmrhQeL7Ccn7pR1m9GjC74r9tqziH5aSxF
uqexFPKINY1jxMLw6Yv5oJomWlbf0cdW/+C7CtZJ5PIvkCd17PZHGCj34He7Xx8VkrK2lTKa0arj
v6qRk0uJQbLaSXbbVhX/L7bbli1vNEssjcw7U3hkJZCw9MKzx3dGkSk02WTq7ZyORY3wNX6XZuTr
pX1jD8+OYNtxwtQrufxFp0ktcdWpqkHTgWfKTBbT57m8NLZRbxa92RKKcNVK0Kq9pM077TU3ROI7
CwDJchzhqeGlZFQH6h3xsd4nG+2y++fkqeXlXVvu2AMAUVmpffh8AY7Qwjg9OttipjkOyx/GLkWe
UxwEU1HduSx/icb4d1LVFgFe8EL8mFRUTuQI/gRL+Ciau/rE+v6zK1B0SWsmhRddcNt7sXrdJjJV
9lT/wmXNCyz/sTIYsr0cBraXGMSwzHODZKbvV8PjFpGq9gFZvPU7WefLfZb3uBmZ9u9aHl+4S288
KXqhUDBBtknULejmWpoY0RJE9IvH9SuLSu27gh+vYPrSXzdI+6R3QuxhDHLEislTEmvJoQ1dzLNN
0aNXDfmUQwHUCEbqWOnkBMRMm5Xr984tsv+b/ogYImhqir/eWosJwgnOJRMpLTP4GhS4HILDs8Iq
xP2HJ5KmVBoJaHxlHIwf/ajK9ufRRniHw08QQgAkEEu8zSATteGw5WssBuMATfltf6w6hS/4L/35
rhuJOVbEYn8rzbz+cdjiyOr0+VGuNjspWQQBPCC1b7lmFOHqOJcu6XryARXbB9K0vEfHBuaPUDtO
Bb9FEJOkDkSBb6n80/XG8jgHT+Migsh6Nr8U5WRNdLD9saMch96xJqEndVPBh4juS/aAF8jt4paj
B/P00tq/YLk1uAZOVt2C5b8Mu/mYasTcPFMO64qXo+dJfL2KpvdIaWynajh06EQMDcZ4Vzh6Bwbw
wIYNeiKVQov0TgGAtB9cCJcrgi5PLBb9m5KD2dQ8ciP13qStiTHfcqC5hnAW5ARVMRHalYwHtSCA
A5BSP07543lfpjug0HRl7sQW3yE5ghgC+ai36YofZ8CXNKurlAROVP5Q2UcNTQRic44OVm1WILs3
8fxN29TcgYNsYKVC/tH/ohoZMod//8eA0KsddaljgVR58eguh2yL9tKrwSNfm6pbEyUEQ5ZhPP4J
cr9zgREIG/ENuYf6dWzG2eKaYj1FueVsoYdHv5EpiQaPqQ25p8mqyJZSdOswLAK0emX6UdDVI23x
xdIubExOpStL+8otDWAuXYPiNXoOuegTFMGs27bngoudBW9Luzj4oByy6UKhsevL44Qcty2VKmYR
0Ku1h1M/dXZ6u3ZJJnnXtbcpcZOauojcH+4ypmw8YfL/5l0L0InPsrzsY9cV6X+SPXqWYBi8vDE+
DrVl0d01is1Mb70N9DT+/S2XMm34XoTTVE+0q8GobERnqS9AzCN7XNJR9JTZTOC/ailNn26EAMQg
ogMQoeZ6DnUP/ZhpfFDUg19nf/2gQJQkfnUS5+FJrZRhI3OT65uPB8vCO4lO/jrA5SOocHsCpqKe
Q7FWZaKNGsNZ5NyX7b+WevZWfDqUkkE8GAlXwChTG5DDH9tVTxTZKjh5bWqMZ2APt8quYPUUG9SW
6nVz4ARD/qnyVMgrgvech0XCfkby3q9+qAy079uDva33IDNxBiGCXvWO7CHoh+h9bBiAZHiWP+Dv
y1vpBSRATXh7Pdlq6jZBGsradPyGu02cbZZbiQHYvibRP7QbUq1HjYbOY5ViZiZDmvBqflMKzuuJ
DEo5PHlbOmzjCoF9LxsLyKRpknyPXkGI4fT0pO6vlDokBPkJ3127ZTYF85P/KbSKJmZUYXdhI0p3
1j+iK+9vDIaorYToLJGSzyeHjbJneMDH9SSmsE/jZlgoBo6s3nwR8OiBBsbeYMYo43tu39zFaxmA
5B0cGLCzHZ1GdPcNvBlqG7Tw3DRdVK2IYOmhLbGMwz96dmZ/dTy9ZQKMM7EAELZo5QEH2R4KNc8q
Cr4gGsm6Qo3ijMha1+h4goHI2KyEojYslWwBjfr7+qXfaguqzi+FfFWMiMk1dRec/JeoUkRBPtYt
aumtwCivudQ7TySoOzWUXm67O+io/4XFLevoqYLhXyIrQV5TODsQ/mJKn09tl28n0wJ+JqhtrGdq
uY6kYLFbY9WsF7UiU4FC8qi8SjbiAlv2wOvmAiIOOkB24mlsvNhFaZZfNVryGbMXi/kraKXOB4A3
wCSZPfr/udjL72Ld39U0kbZ1p50iOA64qTYVvkgNhxi7phokLlLWpfbSNIMGwsM7xSU4g+hhdckT
vJIzn69ke4eeV1p4m4IV4bDCktZvwmqfdUMturnv/OTlOFkpFSk4zAgI3iOQ3ecwZw6OtYAAJW4c
bu1MLPGyArFDNYVEWon2VSLM/dU9LeqVOFhFEWf0UL1jf/I9rvEFz0Cq25MnPkNJsCc5nq+r0d9M
mX5S3Ig+CyOD94l7jPqrgHWgU2qC6E28i5NYmnL7wLnHKy2QA5iuvDIjqZK8j+J5kzvgO7QhOeHb
d2Znt2CsTY/UheBqCqI9SwQBcdq/r7SZyMRwGUrzaRItt7lEKnds3JnPbOmkJHmnNUnNYx9/bDyH
Wym9d2rUYZL3fmQVHCaSuORA97dELt0h4M2DSQVj6DZA6lg0WSHYR5EN2x5P0wLdmD/jsv53Dtik
VtF58BclniV+ofWagNLUQcJj7LHfBA8XDtI/zLogop6kq/X6i0Zu3z/4JFFXbrr3HT8lx9Ny1qRk
bxn6CRb8WSx7YeDGgEDr8qpLHeK+a04F4dSQHhSmwpIwLT76CJ1hE8tvpK6amUJDl9vvsaW+ikso
+oYEyBOaQ1RqMJ0reysmWFJEU8VR0a3aF2z0C5iWTvg/tNOQ7yrCADoX0gDIlrVQTIyLVxfIoTof
YrMuLctbiLSd3cME4fURKBJPzu7cZFN4g9W0dLWrRNaeuJL2f83Ut9KGQ1VBfuIkKtvQwl5m+voU
F5YwxuBIEf9Uog6FPcHoevW4Fg7eoKA3wpQfDopysx5pnUfUvffmbyZ7VCAeLJICoY1xCSpCftDG
zvccVb5cehdAK9jf5sXxOt7mQD50noywFfKjIEZ0My8+oXuoxk68/vtnePw7usMrt4CsLyqb2l9Z
XNVzzLrgZee8zgl97zO15BZrld4SIOqS3saaCf6rvpvZjiyg3OaKb2OaD8VToQoIvpR3FZ2/yUIP
f4TLdy3db/COuZeDIhlaE7qqaU5bkqYBk+tFokpmVnijrt81srHqTpb+2/Rumd+NeNLRONT/A/Xi
bdwh6bZ1WdL9URPh/89U7slBzrkTTJnD1+GutEc8gR5OQasotKZX0fBOXy4dHCa9LKwSBfPO8jbr
m5qNI0n/s6C3KbWQi9t71QxrJkolHHw02NKsXTyLNh+Xpnr3xjN5x0Fun4eMMPZgthqXUJABS0l9
4MLd01Y5ee129tgw4/4EYu7wmzTNcbLLKqznI6SRxIyWmzJZ6tnz8WVbMuu6Z5LJCJAHkmKLzV8N
v1EkaAx+f/gGJAKdzy4ivZZZS1x9+1oibkCu0o0GkWRBnRKrEuG2eevWBLYAn8BSbY91h2iL/7fB
+ddo1tLd2yP9racOWXdoV8x0ukw7JsTQebL52aza3e6F+90AxbLPTnd8feztfksC8/33sTRhuMwo
5EOul/t0Y3JPn6oEhYY8divZ9tUVRPApO4VWMc2+Hr9olpvSmTw879YrLG0YWu34BIW7mc0i+QHh
pLRJneeyBJLJEAOygMndQZmP0IEMl7EXbk3xAMKIqEVxt3AwE2Hw/Md09baJYyFMWOVzLyiyPEd0
M82YyNh9X1oHS1LDFNcC7L5IuV205xedc2X0Pvd7HspQucxcfLs7AIo/QVOcv6Q6fvvGj3e/c7AO
5TR3S5tPxUp4s8u/ZfGmGNRbEAgvY6CQKkYSAJVlglkIhzjPod3oMIlWN3s58uHDRQdOr6uA5o5W
/8RSIcmdpdYYMDJFs9H5RUTYYMEEfv1ar7Q1vAIdQK7RlhPmixM6BHSIM7l4qZd5Mk8zuNc1aM1f
as4iQ0JtLDnxcSrYVd1gLlGStNpWIktJqzJKjiKC7l17txEk9KdP1pW1E/zgcmmBP8HU4p+nuNAD
1Lxdv8OVGrXNFKFUCc28iFg10+ZOLWLC/1YeAnDvSKcRYH5NeOepIuwfpS4crj6lCzwPERrVEfT8
dJL3xdbvUeCZG9AybcwUM/kCNU1tVCgL9r6TPG3IFmSFeMd1x1R1IC+2G+3S5eGJXL8A7TilzTr5
wN3Df9PFiFG/3yTfG8/+E0+JMvGocnyOsuID0S1IQswyv8bON4h7jHEKQZcD/Tsiw6OGVoLVl6W2
oQHRMCK82WM7qZEyMAVs0JzmjgidF0T68GKawmogod2JFLqsUoCTfG0U/tapuxuXpbB7AyKOs9KG
M5ZQfCBIJ4yE9n14W4xRxcK2KLsX+mGd/TG0ym8tHIoNMZItVaiAuTuEu7vZglpXaVT7Z+fkveT2
5hpX6YPvo1ShS9fx+BvUJvPpMTF4iR/TkcFDJqrtzHvuClIjD/9xJkzqfGezf7y7F+Ygz2gqEj8c
ew7QA3D3/+YXFCdKHqRFFVaXHKVKa6GiyDkcLJ63sr0L72aXELaq25NvYOLOXij5pic2HxXZetjW
79yIctt1vGOOpCjGWn/smK3BtgbmqRuA+Npi5J1VnJxy67rwb682JHO0mR+gsS6Y3P4uvmvmVHR2
HkneWN53yrg2KCRgOYCdLtr7ykeEGfPZu3upO2h610H4rmJsY/56m/k5EdHPpi6kCvnO6MnoTNU6
j2GMmIOrYZHIWQdnlt4xPRnY3GoQMrCAIVTQRzvHD9aeeN79+mJW5VwNwGXIdmpjnXa5YH7dcjYz
woR3E00lZzZ+2sit2WYmBwx8aoOlK0nR6vsM6dcS/owunLHjCp0S5gc3hhVeFzXf5rXu0I6MfD3R
nlUZ0pagwOJA5N+M+ORWjtpio6/K9I/i4rWal3j18VFGRPKwsGkvtjYK4IQZu7lO64/peP4xLssO
34F04vCce2Q/BXxgVMY9BdNIE6bDKGXG4zdrx3oPRpKTmmK/t3cDgv9tFnqQeBL+gAY77kha8Fnx
SVRCo5qQHWxRwBXjnvavMmKyV4it4Wba7UBf8cM6afDmf+U3R/Okk98OqFwnz58IJyXPgzRqbAsP
92W8HcLY2AsJfnlOW+NMkKvRBCtvWd0nRSMKtSck6SHBkJggVMFajjH9BeFcfP4vqdKuCQm/6fWO
tjOuV+fKhPjk3AH5Fj9xBI1AQG9vBrY4iryQ0CmAysNYEjPxVjrtNxI9rk5ZppBc6GTPkSLE6x6t
YjG2EKfHiSuvPWizWnp8YZ/uD0mcpyWsIcN2jsSHqiFEFNME4qzpEJZF+9w9f3SHZRKoIKmhxbwq
gtbDx4ZCKyJ6fgbuWWzhubU1gDytZP1yRWJgXFZmGEdPEX9aciBzMD6znOFN0iIuJ3sICbZkqIjK
FVn9pj1Gn7/LoZ6SBf196hc6FwYgsv9ufnZwPgdZ/On6KekS8jOF5qJhwvg/t4EzWgGUGFIFS7lp
sklD6lOA/7kw7D7vid8eP4h3hM+TCVaoCiFUwQ2JZcSPDiHjqjC52sZlpiY/puKzN61gGetW3VK8
EXQxU/NGesWYAmWYOwn9FnL4bpBPwjCWizdHr6q3ld2IQRqplfsubU5QR3CwvJPelOhur/94QO9i
dqf8mTWhq7utX5v3VoBAf9vDlk5Y/eJMMBWkoC+UzAyB0E2pEg35HQMnBld2RpMBuChoWvAWz60l
xG+0tUUlkEA12v1hN1cGzXljaxpBRPSNp7qgEiw6slau3Wb3ySch4bD40TGrp/HK0+euTDo53ath
NouJCUv5zcq67YeVBKU+DuppJhhfYnKSXoiXH1jpEnMYyedqZ6PkL9fpCb29VCDjjhoqz1rzkE7t
/q1bRhZISeWJQ/ord+0ysUUFBxB7SmjuokdduAUt8Bpxw6UhpMWVgzFDxUtm+JivGm50qdJynOyL
tp7NPtHClcSSzw3xJvFwZj5Xx7BSIMZFdcz8iTg0of2c9j2MSiqcL09KrhqKQFRF4WTV8xac12uW
3JT0KU+1mCAdjakoqjy/1lvCiUXHrISE6jdAzGDCDXIPWFaUZrF8qm3MH1mkYXexhkWMcAQTUlYT
26Mhref07PyEff2LAwf1A+0xHjIPOqeo1P1Ipr26JzpvLhbB20fyW9ZugPAEYlF++/u9CnezsK8y
H1x0c5D9cYRs2kZX4kQ/9d56t+Ph1XhkeVu1kbXWje20VPXFpvUUXlfk8LlyRqb0WVMnFgRDJ0dQ
NU2GknWSYYOGnAkaItaS3zYEf9MUbp4t5HQLwsVzoixoPNX3y1TF9UkTGsyb2RAoQ7UAJ+GXGgpr
kzK0+NN01m8hnVVwg1AXL6NvZFFD/9o7z9SM0iZqMG9d8KMTr16AMwIMivmG41mUU/13epcWK600
9+xETSvhxUBx5TqeM2vZpY5nn7Kepe0YQwv8OZqDZKJMrNKZW9Ervsq+Q/1N9z20+A4dLOEFgqJN
KVcQjpe8cw+eHo2OcSUrdb1fu4JFfmHhkebbaTQuL3tpSpST+xSTblcCruThs6D/d87rzFE1vPhP
G1hRJPutqXROAugcVZ604gDDn27+5LaZcmRHVqwgBHm+AM+qBxoh33wAXl8QVd5yRsM9GtMq/Z69
L9oCs+2QcASPNlNqNNOnqHceKkOpK+c58Wmmtj6vJeZHIYNGFl5OPZyuy/A0prXmX05Uk5sU64NQ
DAVcXfjW393lIYjfVVf+s8OZy77OjxQeWM19BV2OBLhqSghBbvY78ATvWVOKAquW4DFIl1nPqauG
vOcGRB+IUq2R3LXeSi+gbZH0D3708BmlWJ3tby5AMZYTU9nciNBpPflVMmBDtQe+ImHzrAKotQKY
375q32PqqdZLvrASEuoWWYFWANk49/9laX7jlj9nDzAgI4zxGvcKTLs042yVAB4ptXosaULTGZSe
xrfsPh/R4iIPHVT8yYQDiDNqeymRt7Ql7t58DP2pwzqjWF3McYN9uQNrhGAC2gy5pvmYmQqLNqlz
vz/cju8+z8GcSwxcSllAeThkzy5FrlVk1T5K0ZOS2P4jDLKLVlLO2mW5epOJtsrYBPRDjU7M8qY+
BnoOU2hB+94Pp9XRbXM44l5cryySYk9J9sNqd3E6kaI3S1aQJiTVIAj3BG+jVJQrrvcO8yBZnwJy
gD9uIqXKI8TugfQPhxmhjqBOnwtIDoh3PntR0Fz/VYDI8rVrtk/W5Kuc2cEPNLKgogLfnXFF+DIE
rrnhLQHlq0V523Xb7pGPrYdO8+Ur5KP9u1MdnXW4kipB3eM4QiJUlLHCY5T6noPhutcUL2qhtBG9
g9j3aSnkm9lIhlMgUfAo63yhpiI2MuBnrEldLfX/HnldJvyyI4LsPR6BM2G9yI0wyAz/lTJu7Xvu
azWJ5be3d14QN5MwVMqK//LvKTE3TC4/l8Lee6lGcvxIY1qJv5IjTQT6kbX2AcZ5GygDMTrYd/zG
fdApOxFzWh4nmt296lhuuWWeAjFuLa9QBZUEeL6HfW18LAQKJJYRRCuzZ050uYVeYhUWgXSG9vg3
DbOJf4/s81AL3HTKh376WJMt8EQMK2/Pg6ong/gpXKr3KslZUAAbYNDf8krGUM57NphN/xhirISJ
hcLmQiiqOMWZaEcgSxdA/uuBOQ685dRY4Cu9y1JfYKsWsSQIccHj27iHjr6AMr+ckHREymHPqAOc
IXDDPrwLGFG1F3DsOLZ0Kugbdk46jOelTTnN0fwExq8ECwPxv0KVfjMv51six+/CqLO8RpbKRGPu
GZ92/X2HWpVR1T4YuRm2I6ouChgBp7hDeQU5amXJd60Yn4ENpeVWYTGCqN3BioqArTfsRRWzyyPZ
gQtp9aPmvRBiEhZwRwEcSUGpP0PrczPhpIHNeQ4uzr08knxuH5mo3bwVA4SycmkLDCBzXbC+Pd6m
dKamAwe3Kj/+rRpUCPI4V0Yn+B8PVqbQvgHxPaFIkYzT7bHgLnPomlotdolXzUGsu4XQIM2krgDS
TQZV/myV7Cljr+V9uofiZ0WCzbOKSFiTQUKWkSzv78QKL2NmZ4mbCklk+vKTkMSDDDEukxo07Ubx
Md4EVZZRGanphLL4ri4AtbzHIr2XDydOo0O+77ry432+1MC2ryqLyggbT/4enzxRdcBqHRZQIQYN
tRkin1/u+djXkJQwufnyxfhHInFuJrqx4Vcwmb8R5E7WOGxrN9y7To+ET79E+uSnoAuUeLsA5xJV
GuuPFr1AW5b7edE5M036nci3TBrxUkat70Ugawu5FEJHu4q3YvIu1OCmp9mKapOdLxwbbVyEElZN
mkFduDKDTTVRMmcc1yC9Bz4igFyj7n0uqRU23AYVQHCmkAXjQjz2lvXACA24A5GkXNFvzUWf8ola
Moydzz/j82YOJYvWYVnWBqmdQYvAbaBB6vdvhtsOqzPL3wxFBdiRioxP062HZcOEe+19qkf2p0UO
FIO50iWQBSlursNO5BpLGPqLaucIa13fY9bwLxWpB1TUAUewC3kJpBqqeopGM1kroSW+xi+6Cr7h
MRLyQIvFximG5d0DJGT4DVshDZ343VERVn4wf5NfrcaYyRLFyiTqStkP+RdH/n1hoqMvpipqOOaN
ro0Oizxe1J/0kiOXhJ4smDuDDSjwNrpLtXNlcEdS08MW/2sGiwD7fmHtbFR2scIacVvVKTUsQOXi
CzPcC+ZhPlYyQR66UuDBoejA7vq+JzzC6xw/EHJZADcU7wX7emV9gqKI+aOyH3/LjwHhwLvSJJcb
IKakJpgKh9JKoMJ1PUrKbbBMocrry99lmdWb8GBmDJ93jdJ2TTXYznNnqlBA/oaLXvRLzuy+ZYaX
wzwiXbNd5LK6eDDTqfHLy8Ml5K4zhtMOqLtxySBg5TtUCM/dWxdGXoD9kqjEDBUhvwjgSroZ17lo
1plYnDcLta+WdFzc456AcU/8lqGq4/gFXfdv3Xl9ThTX+xHPSXW/KUzV3xPp4RJfXNvIpTXfSHJI
7y5yHrxpOtxS5tvS+WnsgYtxWdmkkDEkki21Czmveel8EGjphc3LipAIC8dRKcgGAnrGh+mp9aIm
FgseE2/9AczqhpQ/ETWo/+zNzpMGzGjQB75I98gM4eQkhEXahTf3p28ToLl1Lj3P9R+zrmOdRG3v
s/+2rUQNiajzWMyw8srpeHSrAImD2gK0X/SY1j11Wcvt1EcgVL/GYgZZ2RN6FFsrh0r6ReiHspWG
r+qceSRLFjrfHxh9KVuKZkmS/4zZiZtDzo8ktuYIzZlXlA7bms4pzK+dKGtIizwc+zNWscyB90Zs
IiTt0jjxthD12tkkXMibkDlCV4+IrDaEBSXo+B1dkEy2z7K64hVJjm9Zp9ktTtPMh7roMHtYxsW0
UeeLQTebpzCkNPPxiazkcVSyJc7UAPl20pAkMTAny61sdk/+nQlDb0VFLJwNBJPdR/mUlWkeDpzZ
WaI1uZtgeGvYDml8XBCCvk531NEyMzJtS57k79n92L5vzkM//et3/vqo606cqyZFnsb3hgZlhRoh
ZhFEUeWideRi4hR6rp0Ae8wJ4UcG8aTedfJxhggp7PIlgLdwolcYWTMbiN+ONuLv2ESD4HIWCz7y
+yrr1672kC5itiegIBwhUl/5nLB9EzBCqWxDxEUVYABeYuXFxlMxrLaWxPaEnDqmR+r/hW8uhH5h
rLA7NYDPrE6k7R/rM36MK5sJHu1ovlpPRomBcACq7oOMZXkAre3vliD1frzROvRFJ2rkJ4k2flL+
X4nyEEfQcOW9fEjPxWKoRHygGgs7qtAb5JtwdsDJvx0lAaluWRs+j6hxyqZBhfF39icS/mU+Q6CG
Eh7hXJhxA77GUu9tQq5Z/R81IoAQ5cTvGp4iNXEWn2MKDeIvOUikCuu6sPaVLXgpIE7OYfHv0sKl
Mue9v9UsGxDYOxAww+Wuda8VKHWUItRZejj/5yIzBy0Rz06FlPc30Y4OVMtbeobr3RANyaLLETGy
Qtkzsomj7MkTJiPQL9HB7FeaN5adno9If0KgZW5iypjuWThY6G4UVghEpQm52pkAc1lJ90sAqixc
da3ucygi7/XxSl8amA8sGen+pwa3YG6gmQHqyxxKfyrelYzUhWCDkJtImDm/PhwvryAcH53wijIV
PCwl99msKAQeCj0j7k8RB4QE4vW/E/GI9LkTgjMnpmKdRKOkk4fmH/bg22zMyRE+TTqeH9vjA2Wm
jLk8cD11tanK8vp3PZpX6C8Zp5II5Jjn9ucQldoHO88rcQFcWRwfFJ0FB5hYgGLZnH1d6R/MXvtK
leBbhg6Dg+ylo8l9FbvxmCtzFN+P6ezXOhfKB5uxVLy+CczKxTECLOlw5F+cWMBu41wPyrsrM051
VS9dGTSzrBE269oms+q5nOnLZLFAA1R8DVbx9lNyAXbFhjL/dYMbirBlLeDwaS64/I5ru3D1Lnn5
3iED1XvnZ3SbKED9WRXOiRpn6wbbCKR4VAXZPjPW1ylttcQujh3/gKx9CDtd3zZ4CgwxN+v5tAJt
EGuEEbxt4iiMbgbAVspSl8ULVqPkkjanHr3UR1E6Zd83W8+HQCFnAMLrrHQWgb9cYd/72XGcdpFv
EkZDN8wN0q0iDXgXJrEKMmJryYiaRrV0pepDQSUUBNoyyvyl9sML7UMEicV74LR2XDVnlk/9KQ19
uk44qHQO6tEKqg9X2/zSRmXX+xFGSGHgdurjEOqWYpsDaEtHygztO3OTfx+0uqrnzdNkZr783nU9
hVPRoS2SF4ZATZco0Z4Ru9EJYKf9+P+aTGitLlRb8jtQ+fgDurnmSjdj9WlM7NFAlktNoT9WwALI
/n+y/g7Tv4+4JBef/jVgx1ajxSQFXeGySgGFI+ZrNBj+KcNh0i1PJBmggkrxzOQyUaz5F9yXScof
XcUCNxci9FF4F0ojDY3Ke1fucLaJiRRGwXfCBfnVz56LR32vb05WLsKAlJNqgBTK/mH6FeOsn+vh
4yjeAV+BZb7FlZEzX874M59AMI8IoRU+N0wh1mU9HG1hikIxlWlIPKA5EiGtSu8/vYS6x8J5b5MM
uYqJYToFiyK+ULQaLIelQryUAFd1z9wGlr+ILq2s/BITP/QwsH6XP3dddKuUi/Ts9c9J7D4EmgPR
OiNjlA+BVUrQP0p01Ztrsex3AiG553tM0iZVDrSrayQWQZF8beI7mDCqVkDJml0ViEGH8tUCAsPq
/3wzeeyIF2c0Y9qBRnqnWGKmwnQCKacflLulPbCQXoHgM7JtewVyh3fm5R7wPjz5MKb3KBOPZwb4
btEdDiuRK8pPJ2YvcWEp99AAxO7qdXeP0T1aC0ouIif9YUcrOqf4lrfceFSwQoIRwPg2MZKywslz
A5pe960J1MdD6g172tTbr+V+y/MzibhLuosiIQnRigN27dzC7BBXwjvOEWMweG1k1lqzzjjPJiI7
W/WJm4ion+C/GAhaEcetM+3CaVJ7fgk/1CGYrdYoHChKMPVsIycpzgACuL5UOpv8RLY4XVByupwE
AkLD4VzClzw2tMPjMGNwYRX8iyLBUI3AxKuIs9maC5e0VlyrwORPhqxCC//4u0zQYlspIfotASBd
mNS9Z7zF+oeaHaNfWmB09L94XkqN5vS92TKmQBTyBcEzJL3jpVwlMLFkFjfltRmTfAEUmEma02Sq
Yj+DoUFtmYis3qByeb+MRiSi9dBlWyNOyJVo0DyupoOTvI4INY1XseLnTo3WvBRZf6UXx5H+zXVQ
7oSx526l2KhR9BQsPeW3N6VfFSo1l2XERQXHv1+W/JmBvAVEq/vCASt2oO1KBsU9SF80BaRCo8H3
yGAxTUjEE4efI3etrw92/JpS58zaH7cvN9gxsQEl+F2yw1Ldhf/yuUsTFwqoi8vbkhhLnIyOrv0j
Rs33nwF89gp957APR3qY9cxRIDlxHx38vt57l9BK9tm05d+kMuCu5hGNeMXBe13h1+epEN8xds/a
LOPGUaoFzgaq6X5rzbJFYSOI1ujig0Ke6psk37TQwxL5AVkFlZOjW9CMdQnfMGbHrf+ff7NAoiOM
cJud0d9c0w0vRmxhC74etpw/3/n1JqvFk0vM5jUmfxuRTpzcO8UhZGCEcXkyEUTHOHk1hR1k5HNE
wFWlU9yZ0MBlcw2xkGTLKoz+DOKewqrwU5uS0u10gD8hS30sjJOU5I7AuKyvr3wU228ReqoqV70i
254L3VzA7Jdb62Bqdj4qrmv08/Ms7JdD2/tTElSFPrX0nz/wtu/xfQKioeNHyBtJ5teJiAHWZtHL
WOzRAz/8Y9aX8YAndDt1WGb2rEk1W9sV+R2pYqqbHiG5AwXUEUCDlICZxnQJmE4uWP8hjCujfOkm
acaFlX8R+iEIreDCUdPH+RQwYSuqO3Hc8HvQS5gTOw9s5/viz2oY9eNFFRATUeD0Ihhh0LD2eawi
DVCdftDtazTiwBJxPZyQxhMkS7Zv1Xid7cxdn7UbMxv5yXYFwNpNdnt3RDjlRSlpqj+yzdlno79k
OqNrNyEnSe4sH7GdJBqlfZ1iMviMXkXGXOjivkkyOpC/wE8LShKPTOgr3nLKb57y0CpdLWtTiPOK
0L5W8wAoBK1Xb0JnJlLMz3rk1ldDssqhG+OTztTxfdaRu6msgshbcxQ7P8cECR9/wz7SyeBn3by9
EvrRVaVT2+vfKi1N+Zmpeb7hFxfBe5e81JFaMqqjY77RsZHXINV47WgfKRBtuVmJJ75Y6sCp9AgJ
KEDeLvyO/Qwjv0x+lVTbHxSCcZKdMggc+RTJ1YdRWxxqpWhtO4ms8zjP5yGZPZqoes+/57lWscFY
jJXLYpNjnqkj4n3fDwDVG5YHMPlLM9Sft0IvpviMiGos4bl9oI/2iTEzGpginDUW/jF43f9w/LrS
kKsU3lfTcrrSPRdvGZJhvCK7kzmxt3mADjJ28ncOB0hQpRQ/88SC8aO09UR/P0RyYGdA4HvMQVI+
aWYRl5NrvOhvjkZlDDDf3BjT9h2yb9Bqv5lO8j1+jf2DQg5O/zkwyRn830oV/xZIn/fbGFQx/I1a
MsK9bbepu5GNDU/v4PTuFpuJ3pdY+6hiBAR2Go3QYglY7qU6kequ0BeINNdrgbcl4vfTBkfZubQy
Gk3D3VnmdhFKULpe5g+OSaf6MPHcx09SEAbRUCDfOFIm6a/aDUOy8ePa1kDFEna3Rs2Q5vvJ6E69
aBEaPmakqp7gYZVLvHX+5Ai30/crrqjv3huR0550eWHLWDtyPrD0jC2olPWBM8CMIedOcKoREq/B
34K3R8q+sbIUid/8C159VnF3jlDg12omVf864NnMePV2maQSdRsVXpdiNiQlcVVk9wu5/SMEGOeB
hXi7bTDnmoXYZe6gOwthk0SYFQAtIo342b2ySKwSfNkciXUmulXE2ep2oeSGoPw6fhsn7im8PvQl
8KeC/YP0Mf+GvCPtoS7/wH9+82tG0gXT4YODO0ZWKu7i4WRPoBvAZPfJ3QIDstyz/i1f0VH4cj5W
0CjoDWMCW5mDKsal/hJudABxd5uWxeIJgnvJWzoja4mUGYqXTOI3NaInod+gA9KNwVnvNjqPdhTv
tbKFTPESlH0nOL+8DS0BX02P4jvKgnPNBHHVc8IBg0sUYlKrXxegwZeSccpA+59b8JoY68ROY7Ot
Y67+EwFi7OrUNk8JpRtJNbnGBV8ej7+q5C22hLZgmQAK3Z4LTUKvxtj2zvF/nH39PCftnvzymt4m
sFN76bJ1RaUIgPzFzXmkbTdy5cETjFDtdcY9ylfEDCU72nC5dp9KT2nRjLfl3us6ke6ZKOe11mGt
D8xi2zG9M1g4j/8PMFYW5kRLzAkDi2CGk01JSLtXQdMJRE7Tjd0yym9R9kul5bxEcadGFCwo7Pye
ww1GlmgLSMdI8bzN84P9TIRg0qwU/tQoThqFY4lBxfnFYNAvMsU0ZX2D2IbchRTrMoM+Gzib9kXj
AwYQi4dYy5QkRNLsy4oZNSWRjEwC4enfCYamkcuoJhToFTnCB8N9deKrgJWvpako2KGnWvNSBDqK
iQkPV/e+jFZ+gOiWdcxTqwoPZrdhcqJM1JgleItW7O0yaJki7QkNzic+/xXjYuQiENdQJMUTpWGD
+Jb10oxOjAQTkqmmL2vrBrs5x6Xk8gxqiZDgVVYIRK0ffdTm9ZKLAZd+WjXNLpzbC2Jn8s3yll6h
qpfnLVat8KBpN0jCpBElDi9iJPAUI6SpIiM8Ei8lUYM3uZnKsuJNOMsl0roA/+UtSa+/fHXeyUO5
qDotRf/INgpn9JIOGtoZ//5OVGpnV9n4wecJS8JcyBZiZltSWF1pXe/VhwcB5+nzJexxlwUmNea/
7fMsoT9Ce86i+UcB7BIFr7g6jBfLg3tNYrSjZLr/06qTKqhpRYi1K4O63PKYv/4Ccc8GL0jgnfpP
gYkl0aFrZN77WmcrIAkPEP4tBiueluwYumJ1X+2D08Xxa/LzG5zY52L8JHWz5a7y/4edDBYVokAW
qQ92LvUtiFZMILTg4F0LKbE1hpGi9WAEbS0/tjHFgJ3hZky6Qwb8aKVdDmG2tBCaWBCnAeDpbAY9
8ozuSzopSr0FN3scuxgrka7k2OCQH9OR3I3e26fauGaFeNuCwPmoo8Ga1FvC6n+GtybQG27qgW17
FXYXjoL3rpA4J5MlBqNhtQBO8r8uUiOqiU6FeghI2/cxGzc4oVh/vLqmQz94GVPLPF6bickK3GdH
1HrEPDQCugyPj8wTCCJMMfSphy6Oto5GaLdAPXSvewMqGyA3j6Xk/nlghZ1ZwTumWij+Qm8QViAS
rIbhJl83B8/Yd2abGTiD8sgGjI0o86zhca9F9xGTSOOr3tr1q8+nhGkWZqfCsgiqBhRaQggHSKml
JCENZ3O2dRHAU7Ut6b1AWzYnokbwleuW48Iwra3eYJjJmgXRWBvqoxBYOM3FsCvKvVwaBNgzoOBx
TZjebQkvSgFDKiY+XMiT5eGClyjY5fWQn33fuEEdEX3bZC9aTzUXzCuPWgj9NjU4lUcYtpwJljyZ
GNOx/9JdnCFa0WC7HsXY0R4F0gs1hIW3icjwyz/bFKO4qD63fYa3TPAvZF9N4oYuPwxyD3WyBXMo
G7M3cPjFwMuiily0MofME+VDW9qeQ8D71DOwMiWzx7Jzccu9xzpd4dlBfNFJySqad22S61TWHhfC
e3k43N8YmqKnVVfvQPGfihg1t2Ti22E81vNiorY0mjhSshZ0ZvJ4BBV4w2NbEafmHcg4C0SfWnIP
qLTud1wXTvk5EXRhcEstqoFQH+XCOKEklBWE/x1/uKWzYvkjfkccx82vkL3bbLuz3tnCK4A/lSmo
Iz3uD7PG8lXYs5ipIa0DooUy2eDf416AD0+rcqYGi36BBYnxylWcwOJxzd21Vnh7XmVejnBJPzj4
odrzqHDEqnq6RQeW3iV0x7MmBkU26mNWZSGkqxrIj4eyQWIjNXWd9VlkOBMMhfTaNOHuRvX35JYu
d1mI6I0OYgSHBVwR6zjg8FpZRGYcFMTSsqP+t2aNqdClL7Y8j68+Un/Kzoz1bBV58Va9rF3t3mOU
sFwjxJYvjp5+f48GEWIWzQEwIheqjVrh0RlTafxRf930YaqlS6VgUFpg50l5+GexqDg3hLmRz8K3
zoMIRyW81o9FbIPXHbOWhp2O+LNdKf4aq7aqq4fT3IkSjonKrKxNWfELyVJkjLM10NboSvplX78d
PMS4HCZCXCFwv1EkfmzGZW7zwxdjRStfZzBfHeQ4paCjIcOlAbwg+KbuX1GhgsyggZyuAQABa5TH
o13nouHF2qbrcehNMBFwY8PEYqrp3158d6k5YoSTaL5PY8GZd/LAbLngsu+nVSdvPzeXj3qkRrjp
1SsbNXANT23rk3ZiPY7aZHVXDwz7KajhyEWAkIM20gKFggZxrPkuEmt9uR/ewP7bon9hXLCx0K91
slErko0yVAyGnN/SGANUvO218QqXDircSQn6sgyu0A/d3oc7sRSFnkyLxwewq9GevYnntzzcOXz/
9KMxLduOUCUKB2tDf7ZocoA7xwazyOYa3/0rVnHQDMEtS/UQ6exX1iVbqRH+aD63oSFLVwQPu8Ji
1GilLA+eLIa+3tjGV9ZgIX+95upOcTEobF9GtiZ/94YCfGsaMjhvrys+wDEOExmO1t8P4dE+uyt7
76DHTKeZtyTmSqKhTENeTLkftlJFuHEiGa4/+rNuv8Xu805masm8gZseg7s4e5FpUVnZea1NdRE9
bLc/53xHXLqHGdMpYDDdczvsf5virj/xh8uv7ahOW5U0Ovz15VpNT7gRUJCfWridDLOW5sungzxh
rMV2f7MtkR4vdEAgcF4XN/b5THBNmFG845HqoCgNnp1sqSQL5JlpbPmw4AmZeSs39eRhwT31Wfep
xPcjZpZTbmTe5nBfF8FrOQsyNQlX571Vz/XeC9I2cm14qwqC4kK1M969Ia0+erIYHjgZ3kpofOUN
R1ldNiISzTo6vpE669z1QUXEqyeJ51TWGb6p+bMOkqUQQnFxFb+gjCBcDA8iL/4/F3FhpeZCxsrf
a/5FAQjbucS8eN2fkqOwxQD/6v28yd6KTfHR8iE+RsAbuPFKSstsNxm3hppN4zpEDZdx7Ri6YIZC
YaXmTd3hNQhn+Be/UriOQY2TKb17KH+wD0laT5VPx10LaBgVk8hbWgCbehSUZhcIHA/gSxqFsX2r
RzwIQuepcKLVsJP+VPQC53ER/qokCmTGQKKn5MkzkIzojm8gsz6Ib+k5qM8YZKxJjnMPK2UBE7eA
JxnbycLKDU8p9nrUrcgganKgCr7YdKDtpT3QIOcZ0rDSYyQxsQb3xZqFX3vmexzBXma2xDMttVMb
IMtXTiW6EUKOBQD9V5MYJO8iQ/L3G04sFEdo56DatdlboL9AAPfW6wW9IeYd0xz9tvmGAzeDrrZv
1aJgHHO2/aAaz6Arm41/VNehabEGxUXbLi7ejSt2CgNdBFrYW5hP58g26vODTLsFs+iH83tFeZUd
XY4j1GUwdL6YAn8Jb/l6fO1x/nQtPkBFEISynLe6CctkI+4+4Kjw8G9Ug/YQVW/khRcS6ZGPBfrk
XUQ48wumNTHFJYpMn43FukgaizGYuDP9KokdeEEKoS8PUzbAlPXw7o9o1ovjSS0N4zd8woflah15
RATHLZgWUWwnvF6CsgtiJwuhc7dHopMV+JNis5Xo9iHlz4KmJrxYOTm2pyUcEOJss8yfi89UBR9G
6lLkArt4ySNdVIQYMv34t6G4ERrb6KvvIZJKA79LyjywtarI7VUEGw9MPy1BZSrC2EDqI+3S9zxO
xXsuubPWcv+nWqogZRRS5VDnx4yXtPVbZCIEEIqug4JB/0jIvETj5rBwpg06R0SkE3O67xaGYJzT
InM1LiE+7tkVPxAz9fxPPWEb1JNjjKqzGwQS7TwfBMKOM0yXF2xtIg02PZP/jqnxnl1fa5FHSZCS
aYczFYubqmQPX4mEptGGtxGkyM8QOWH1msQ7MxQU6kWvmumLoM1EuAwcPG/oFVgEdivg4Jd+9J6P
iRMU6QW0g+2SIVTjIxPoThEX8IU6rJkurnflgIYlGLP/TG3x0h31kHklkqi/237D1ihMYJ/ZX5mE
C6ygqa70qCEtlTJSYWMbicf6+ih5rHc+sENFTwwjIjyjtqVCgGz/Q3jjvfmI0r6mnU47mCB6Y4JW
8ysEvjXhwkPibF2MMSbFBTeGOtvNQjMJzQeidzo1XZOiZqiUdef1Yevla6wD/pm2D3I9HWk6d8UW
TbEjrzNKuNjzYyPQTvALJQESb6azTyfdyKsv2yYJBFjlczoirlzon6JdBKKkm2VAVNz1Y3XGqeDb
V8xPsFanv8fT6U7rBcs+G89bK93bIOMO4Lhq4MICic5vlbdEfP1zU9Lmjf4eTCYvkMmaevwpg/gk
KpM+hWFEJ+AVNXdfTyGXT1xYbRCzRfRn7iRa+Pj+fL9CFvlAlhwMyzfOXQcvhqDm4EHJBcDZ6JNa
PADjqG58xB2zVpWRnGH/fk+iW+nMt9cAZjyUtxWFe84Ni5qkE/W22rqam60vXTaPWisdey74HtG+
dsgmkTlKKfsLNr283IFkZjAdYJhEwya6/3OSUS/b82TnuFsKCKFwRLhdsg5p4+7jzZgIjfCnLidJ
lV1eRODGjC8jpmkezGlHn87XM1HzRJViQzzq7suoMYgagApKyYqIc+c/e343GwqfaMySnbCWvVcm
C1bI4cHMD/QG8VR9dLRDsAJL9TdR5X0zxUycsTDEA7rBiQm/4eErqLiq45Py+0CHNo1ZG56VgKPQ
cjaJaY2qXZv8osgVm4nNrwxTDwIhc105uHvQqABtbvh75vT7EPy3iO4hm/lCRvIA+kjSvnn4tDO+
GsEgjd8mKmPzOyeVncqtMl5ljCirIeaHI56j51OnsSaNuNa4RpnyzdleB0nbukQHj0VGbsb9cGx6
JxLhTkLS8f5Ow+urfyEyTrf8I1k32cewT+UkEwC4zcMhN5o5GBrcZd4ymRMVjWXZHhoWcWRb5b/R
y74oSorzi8KBN1tE1Zh1Aretstb3YuP7/N/E1vQyEHUWgbSrJBk79fyrbu9gi5tPFfTwaXG/kH+y
MIV0KN/6hd0BvGIOCLG2YLKxqMG8Xr278NiA3vYiuj9iC4hZpAW5qIEjwVZX0+7vrEktxv0ltQgs
jZiRewjxq9DdyKfMF8JEs2wPpI4nSSC93czC2bO8Dc57Jvp5QGbaByLIZ7k9309qEgetuDAV5qe9
8WI3OweCU7ghrGnu3OvKCtFZiBU1FR5HX4CcMTI34u3MmF+X68fh7ppCgv405U9oIByYryvT2qXw
uh+G2gSZrgW3bswwbgbegRU5wv3vG/fVRhUe7HM2Ft8KqjBXQ6kkVEmIIPKYBQxgEDWK1t1K3iQV
4MykUiaNF1zsvt/JsHntNaqbHTQ+Z611YIQT984NZba0X4dQkfHakEuqJdsBhu5qHIy7ynxtrVv+
kHdJcFSgRbw2uISfd2SfU6TyKDnDZEOf9Lji8+1jU8h7zf1dVozWfYEl8vjWDXPJYPXDLbR1nKi4
Cp6nqAjpGVuRjQkSw4INjUcaf+wB0mbL0uLd1mDx3OJy06f7L6L6vLXRIgT8oW7oCB1P/6OO6gS1
yQ4KEskHCcFUMagc/XWVLiGCOZf4WJZaKpbxO1VL88dE8iFi4QnIu3314LcKAU0jq6GSfb8VFwNb
36l9qZVZIMma/56M7CH+37e9LUju84aCzwOfJMV3MMRInuoZ3kgm+I6XWaZklB6g2U8SHG/3Bi9L
AS04PaqqJ74CthUlWKoX0oQvPh86ddj1IamX/ZzGe+XET9XGbUe/AJu6doH/7VbgD1hin99NlnSz
I2F3kS67KngY9Pu4fcd3Xe1MTjrvzrkAzNT1WgH27WAnuaufZ3KjLZRv7IEduGGO/rxaFGDomInl
GL0merR9lYEm3DqyMAuo63s1fDWCqN1id3PaJ1YjodyW2SxfZEJiv6v0US27a8zVEfxK0fExDvnb
sPXoayEnqUARv5g+dJmipVq/dsu8HJ32U+Jh38nn4ACqMTyVPaq/OpvCEMJOMHg2SmCt0G+ty0Nc
E4tTQ+jidMB5I4sxGo+XOTIO+1kptJIGxactMIATTdqQxUXUYCN0YMCkxkzUAbqWc5wYt4v4+dOd
j41ap5idzSJlgGQAZ4FEi+gxYqFX7hCggO7FLBUTlUTp3QHPvMTz1Luyj1216jWAQsqnuxh/kZxJ
a/2WLThg1LanY3nvZ/eSmRIxXNoewIwrcVfiDAMsucUrHRdRRNYkKhGPnuf04kOliCGcwcbJhJrQ
1AU/cNY6iacPst7xPJF9hYeyB0ugQMkKYBEvI1y+DvmuRtABqpGXFPYJLELxfpJmxqUqWhKw120Q
69eV1wCIsr47D1fcLXTZk/Xtq7Wf4cK5wPbukW73LmAcCTFguVK0z44alzr2nYwu2EcynC9TAxlY
GaR1QDDW5bk1zHq6W7rQlX0Ta2eWA1SIi8jQ/W5AKdThLiXn5AR90Jlp2nRowQRyzYS18y1MOjpV
UMtLTNXy7l7tX44IeK7hZBU7wwVBXYY/vD4EZZ2x/3LxNxGLCSsQHWSqzFavhRyj+5Su6GR4ElNN
ryqtB9wDOjaKAupYw6dDgn+wJzCEZTkBOQQsphwoo5UsK3KmMpHM4ovfxlAT1qyjSZf5s+f8oM/Q
b2YChyc6ljaGBqzu6O6tKBhiYWcYSkhUMA+XAjAdF9y2PX5wk8ufoFZxoNI6i4mep60sSh5s2i8J
8fDTuaBz8Xgtqv8Y8WA8xTMKgKsWkftJM9HXzablJiT18Dz5nXunYeqBSbzW0ByTDZrH57O28LCz
e9Ghl/Ep7jOK/zeca1Yzh2yr06RBUCCszibssO2MbPeLDLsWma4kJ23AqkB3EQ/tR7wtfmFmpN+v
QP/YzOWwHerfbhdrJ+Fz3I/oq+KIxw0Y/kbVFWOKNQhIjWBS/xE4d3Gqd141jis4Ue67uFnuMmHP
m0X5Wp3lhvhCd1VwO5tlaTCo2wsH9aAEtdTfFnQVw5SAm1r9+Mhsnck9lPKK2o7TL04psf16gq5X
r8JcBG4OT3sebsoWfjrLX3G1vm77+tR4IvjID2LXV06eIq6FHjdgaGjqFMVisEkMbIP0sjh8sMzO
Poj43+STqNoo3uyYo7kiKFEsmT1tsWdA0mGCJ4SR/qLG4OE0diph18lunQ9GZtLfJebhlpLnig+7
uHxASX5qbV2Zv6Oy22fT0U6E+H6HRstPGwT+A+eBvNU03z29cZvYCHGySMmGbbsKfjn7GMT3fWjc
6iwFgWUL4xbyOTWQAu1oO3mG862MXdFsRT1NwcR8kCTjvQ4m8b5tK313UEigCiDcx5EbIkEzfMCy
ZIMwa3lWRndiyZfS2cjXo+pKmM8alt5kzGWCiYPHf4UBpEV5QDdU9Ov3rBWDAmiGIlOT9oyGUUdU
pgCJenWNR9+bEjpgHLWAuO28CnxtUJucFS2/M2yqx4IZ8P4R3BGB6gRCf6sb50pl15O5pJa2RYiF
QKdtrFO91OXW/sADcmfWSykT1totpIPjy+peKVQjhSFJMRuVzfDViNJol7cVTIyowOjmPPL8E2Dc
btVgpiAJFjBBMtJAzj8MA49HIdQdeQ2Qa7vazZoBKhsj6m7ktfj2UTK6kyRzEv23GpggZ2q9lk2L
qZSajAKZxeyz1n+3/7L3zrdtxOZI56gw3qVW3eGwX3q3yarciIFWNaawd45ix7H6m2CxO8jk3yTJ
MTR6I4AY5dKj12a7ibcmvAdz4PEvztLW3l4rFWrYFScOXmDlvfKTfDRRtaWU4EWSdtjS++SLrpu3
QwNITZzmVObCKThDHrCdC/FPC1uED3DYs/JIykAE/a1KhaatVjK4oAxQhnIXp4nj9o8dDEzT2adH
e4y6LrIL87TggrpJRn0TqKila8fnWzgCswheqjIsnVATm0XCJErNJ1oCfuGMYCfl/X0IQqV2dzU0
Ec+DfTdE+7arITbpwFu19UKQZmIwMScyRQtjR85sW1NUb9aRCCHiIqkIcWt3xynWgc2jRB3uXEUi
9GxPOOXnbUCkcZEF5EnbMIFkjY/RdQG51ZaygQb4BLYKi+nDxXOxF6FuNn+3wkvPzWfCvMBmQ3sn
xwecsiPYYPSGYx6yJCozGEbHuVnd+0abbA6+EK4953FV7ewMkwcQqXNJbk1A2soV5S2iyfoKp7tk
kWnZf/Q3X3wmfM5mKifi9BCyfk8EmzueXCd2AwIWcHvxk7kRcLW8ET3lIAPI2o7sFjMrajD2Pl0r
AWdBdx4UH09in0M/D7f0ujN6euaMfxjYcUerhJMkwF3LzAvhkEv8JQcHPH7s3bKUkahGZ7cMLNq5
gJ93nsoDL8Y6rMEGkXY6vrCwEfSAZosH82q8pCqMsdB6fSZlll/LAWSewEh2YJlxsedkWoC/MdW6
E/u+HiMu8Zt4mzKWFKQvAG0y2FuoJs1cymHqGgii/MuPNxHOTXUmyoxSH6Xgyc7fiODBU+lyuOd7
84buCnTG7FIXZBdKY5o20FFkFqYiEmJUIqYQh68gGC3WVftorlxU8dVPkyBcgZ9+PCGqSbg8ialN
QF/A/pNSW81vmi8j0fr3R2qTX4B/5zqY63edb/QT0i22tTt5pNfjvkcKAZF+MQ/9CDG07xCoghIH
4LuHyXjAmvmVhugFB5K1kuOUzZ2F5wHltnFANv0pPyDv+AAXHSylg7ml8UKITdqZCA0em+JiXmg+
cLnYgatNkehpZk3qGorI4Zo1pxM3u5J8btyPkZwQksJGu+SoBTXDs/ZX1M6tgHtXPqHISoa6ANBt
ZWfGNrs05eKHspJY/1QmH8ath5LrhruW0Cb/fyaIvGkRPO/2XfZBzCKNMWwAUoVXsZtAaNtYLQa1
DuaixBhc9gX6mDZRJ1YovX6LjUihl2mOUCWZhx9iDNYQ/JPptI67oe+rzbmXqb975v+ToLbKeqbM
llZ002VgpSdcFl1JXrJV5TyNrUiXBuPIYd4CAbVphZqxWGTgaQXZNQK8w+wyZIk1spA2Y2GBOk+P
+3pFmdEfZaak96DhKlIBiZTUQoa73vS6IGCyigkf674gV/tLOr4ry6wKC5tZmzP9de10IpMw/ugi
gU3gzBNE+BgVCsB1JOyrVBUEsFElRyaQ7uG8AbirKqEv+gy59DzlHUAPpNJB/4MuE1j2ZITykfxb
AqA1bvg/7CaXxrkm+oMLMpckdmvbPb7bK+bgQmgQMHMirn2NZh0AoLtwyTi/zkOoliGPud7semV8
JM+rvvKtJ6oftYQovcpz9Kc5Ga/N/rXToQ2zeW71yuXJ0fUG3BkmY3NmoW/eaxezguulKCaRbvXM
OF26X48gY+Y+fd+30NsPUbzGeNayIJUKonaaYUv59XcnpBME/LJyKdLW1Jb+jAQAbdMikaU+Hn2F
C1nMqot04H8DfD+a2hwIMkplbpcF4qAbdw9eDRX39OC0IvF2rVQV+iKWuQHtPK/1nf0fwR6NjTnE
5ilv7Fzg7vUAO/VjXU5tLJqiyVBCPCZtVFAowIfr0klJ9mUW/0B6UkFwpe3oW7li1o5Km/8A6ZHL
grSeu9A4aDXhElCriASWiGMHGp3bmPUd9Ap6N9XrbYN/JNTI2b6Vjaucmgi0b31G2KJrQku6/0q7
vsXD6c+wZqtSrvdccqatpqdLH+K3i/n3ePfLv7OZAOKEJCMYh4PFjJRypBYyHrP8eQw9BqWCFpo0
DTFHHtKP30bziW20aGlQAmVf+7BIJQ4whDCuVO5POHKz+wVJsxLpKzwPEA5RYloACgubHLQcHwLw
MgewK6P9Uh6kFT0qGsCYDYQ4y05QNmdpfpghdmUXJecl0y5bI0vhOMjv9qdZY8RWQegZzNrrRGRs
o5jvL1a122+21skDXXP3mjCZe1/W1Ps+EOIrArt9wCZtGNzG5EVv4eKst8NqdirqLvKknBgqUApT
OdkEUb97juHOpgRtPY9SxjcthXVjsT71QiCQFtDEBO6Ni9RvuAmc9F8QEW/S4MaPr8S5VbF4gUP3
2ZBDuNUlBx5Tt0zEVkdceyMwBeILj5xytW91KQHpFLUaYCgQbYGgMIDJPAKOyRT7dgYnB2ksT0iY
iHoOJo6ahmZK63DFF4R1CJAw7rlLl90CciiEe5D0H9b8bA7Xea4cPIUg2mOLr85TDAjTJdzAGApj
l75OYGdAy6Y5ahXu1wrmLA1RNvWYACE9GcfwYvvHZnu30Kize0IOIJtTlYVUfrsDq7Aq11an/Ydh
NtaRSRnZukNfYlpeBnMU3R+y0chbHtkq5AspOBN+F6yBLIvIqf5gNIxwVOGWCp4scGLaCmA0lCM4
unUoXMhFXe/fNt++fWAj+hT5xJxw80mNzre5INL6fxf0g5Hn3wlnu6ruf/IcFUPdleCNZlhglESE
pjEVRGamLBIf8VVIjXvfJi+T5vMqjzzRK1xPhyGpVvMm9LjiF0/NEG2RUhWR+Srwq2zDTYDHHRKx
upLHCBGktypZg+K4ccfXqSN+VfvGMXf04gzsymH/MOAfN0adAIDzhaB6RL3OEcsZaSUdT6sk/RA/
GdofkeF6zobDM4l2AKjnyVD/4Qttj9APr5gS5+UZRnMTMlxV8WVkuiFUFjfaGRgYgmJmrAco4x+w
bMJ7mLrIK2o9jSqKrUuVLJwfDDcDoEd//QymdCPwUWqaIlGMD1T07pwKD7+YnPII7CiSp4CD4Gs7
bm9QAbyMhbshQBxQEoNMwOTaYeLRMN1yJ7CUfx3Lav580cilyC9VD3KogU01mwwZWgvi4StUBwV3
A8xRMsxtY+UD8Q37zBY73OYZoo3rPHuaPqV4i48bUPDhXjV0q0qDpVw8IqKUJ1SZ8LyhXsIw2A2g
GfptSK9FQf5dBxEUrR6aK3ibiY47vzxqzanYkgOVBzPCWNu6AJCcNROsSDa90XfWrkzEXW5oZJK2
0axwaqQRTtMyTqEkFnRBtTblV12nHkWEzk9H+Hzi5RBOAqogT2JeiNnI7Y3MfyYcdWdtGmmu7bKI
hvEbrCdB7Gcqh41SQZnJxw4sJ8UZPZ78vB1fE6OXVsQ/YbHFavZmKy4adpmuRLV/ovYgX6Mi5+oX
HqI1zhI3XdRQZXMyeG3zOfVChGdvqUuwluzPfGw8ibWU/0vpvz+ghqt9ypjW6eZMsj6XXPO4JbUC
QQBSa9mkjH1PWDn+ge/DoeEI9gurcC3hKl5dhOEsLSZOvikQKCjMT1JpFIfsVST99zxM+KQwmF5h
dWJGqMc68c13qF9pP4o79q8zrv6WVBksv2PsLB0Yo2D3uuxpOk4fcOseWQ841W45xKLk9MtESiSV
2pNJ0BO0XonCOtTbEUVQHBvzJh3ssndnt3lqDeSV7bn8+btEiCXvAz8xAV/tLbUhb2LUKJspLvla
zwX9JMUk4cKf0VsQLlgpBnr39pA+U4bOs60Kov5ztM3T2nR45iQQ6w+To92x9N1SViJ2VXnTvZFD
v9ShnHRJBUkzKhNbcnwXnsaFwf5YbST2TtUlE8r2wR2EwNGgd7Ux+8etp6iOXUM2QXqxsdr/OnJI
MbjyExodxpmu+WzvwPZET0TawMwVsSAkEkWMxzysRgY0LkV42lGJMbiVFDcDi7VLTAgaNzWEoC43
iLwMACGiNLcLZLIDoA23t4BWWlLE+ZTVjK3XvLzQzBgXbNrLwfkoDx9ptwskCd69RbP7bCMUR7/6
EWw/YlmAgy7keM4C5MsfhRhJFjysJPhnaz2R1HMFmk7lGLHyqDxN+Rz9gtCuyPBDFE1SX3rJpt+J
tilvpeLjPPSfMiHJo7fGwonzb8JYJgGTPKn4hlMNOpw+D0fMGHCXGfEyK2xYoI8d9bO0G1F5V8+S
5WEpWsLUXW2cJHP2TC/XLUUcju/n1txiXrZTMShspmK5YqbqMk1ZEtDEBiO5vSADrtiPbdqCPSyz
RPoFRFGLtmKdnwPiFYRic4vqDS6xu1i0KbEEDSkFy84GM39r5lsNinka2CPDP+xrKzB8q1MI6NoI
B77+PS7zDGoq6FSnGAlfrJ9LKcJzT5lU6nZqiaY7lhwYYiRek93l2jva2PnCSjp+DKjMl/v58+Oa
mwBpabCrOFHoaGwFrF4mTaqS0qqz1wHePe+GixUdb4p60OyWC1RcEVgtdCzkO+nNmXY0O5LIfp4Z
YSJeWNgbWYT6TCNJ/3l/D7y8WtTbn4G9cjj00TbMdn7EN7TJpd78i1s6f+IJ5ahRsB+7+XsdVHiT
LAQb4xK20WZnhIsujdtuyjVEa6sSB36hT+n8fGh/loIhSDEoiktt7YrkFChoSLfYrKFdR9KtPayp
SjJAFlgJQbnzok4QEZPiBTPnFxG1ulhbCykcOGYbD35E4RSzrvFZPcuywZwPo2/GBH4FxlTD4s9D
QrRrQ6pRESsfzBumUPeEbR3csB5NZVwNP/04DWq6hNUR4LTwX772Ia5NzWkyQggUd5lPI7raxsmR
NMb93X9WRkClS2L7NsDURRBmg0gM8SNmW2Kf0NTJ6Y5vPLWPY7sy1dWwqG8SzPStiD8qL8oZ4zzT
5sCeJQnWtiRpeSF+kw0K4KQovIZGUX7J52dE2bbtnmrzP0lwktRA7ulUpyRQ+nsL+UynbLmmkjpm
Ps501Ezxn9Oldi26du8zXZMDU8pZUg4d9f8HpVGQrAiNG7+OfvwtJx4oF0pI47dY0nsjA9VI4eyO
pFPaf2Qp0FQfqYOEJGU4YXXR6thglK2fwhRwOh8VZ1qmk03k3xB1WJXpSjAy5NMvSlfWJgpHdG9m
dirVNv3mLWJr9eqN8QSg4DNDgs0vQoSIqOrcHe4iecuct49jAySsJpDnnuDmnBRcYAL7BiDB+o7l
0tTpWHl0mgpyjbWLI3OieEnWtR8lH4inRe/RLvaoPY0SfXFYHeq2v5bdx3LX8fFpwd7Jpi8aTRaD
27dmXiBIHxkQfgUwVHM+YgCgotHSNh+SAQUhJVIeNzSi7lV/ouF6ZmPPVvJ182sKncXhJB4oalxm
l1kvA2VRbLhukNToLKmyE16+LlYhKUQ4PQcqj5ahmJD90YjmeyGF6++aAIaSdoFoHdWCAYXp325U
mW0maDFxdeQpqVsSIvWaGEqD+3uXJ6cQ0vyBTE91ToxihUZ9emxCPBM43GKrik5UAudYHb6neGNd
ZRSyM9Wg+BJAZXrCijn6uK3HV9VOslbSbUdbHOPj5mRZddBPTUZ65kotr/z3VAeyRDgEpSeOHhhH
9YKdFiKBWrdwO68uRr7MtfixgMqbY3SZLfxFT3JIFJEIyWHsyoGqk/yL7R8nXnfiXPYmF7bAaCst
B9jLA/UjUPYF9owI5aCoX+Zx4ZGHjfSEQ9KSuOeTjxlXO+Ova4ma9qFoMj4pqPfn4Uk1j6K2RmgJ
RZKsY9kilSpAUkT8SzYHfJ06U2dzo3XgRIvrTM1P7YZCh+0DqqAlEKU5X9OrVqfFegnJjJDlfXMT
XpmmeBQzG/r/xZJyvec+1CK5l3/PVGW742eKNZhrrlHSt/tbIyqkM2wh7n8BbS5nnh2l6Ia7qdZW
t4HMuMRoShMWfKoGUq0bDyWirczqs4GeK/OKRoulIn6LinpV73M2JMo6PSP16OvPGjvcDAY3V/7K
oRzuchIRMc0zywCg2MB+l1QD816Bhkzm+K4zjW9Oz8WZRrO7zjG1i5LIWWN9zlQ98xBIFlR6bL73
SrTCmQ+ywn+6/IV9mVrv9gQL+X8v3/iiDC4n4BJncAA4KSO59Og2RC6oIV8vNzEP7F/Urt1Jnvtc
dbn/Bn47c8ogicYeS2IpdSZRAm692ejIryk4IWqEC3gBvXEzZzNF9SpCaKxZ+1tCqVRPll7acW+F
SMrFLdjyVAk2dyeDHF/oi1HI9LkwTiz4jA8Z/f8TFAmK1zLAjx7mEjpusZAwXNnwc1cEdLOvHoR6
EIXHAWd0Wjif1UL9bHTF8xGAUGAxF2HQhiaVZZmqYVappYGmj7PhVM9KBBUKmYyy2o/bHXfMIRQn
95qsPW/U5conjgSL86lodFAqEy7eFfmS0k/9qwXXl4/Tj6Mzqi0zRFacTa/Bar1nTIx0Ei+az5Vr
qNU2vJcaRvFpPv+4kjzv+I1s8bfj/fDnMkWGgSG+b4JjgAmrfbXnx6uhkqTXYaBpQpBSkfpqE/kl
b8z1Mwv8S7FcGFxc5suZWTq4Rj2UzX6EsQGjof4UgD03s6jtkKgPdpDnEP3RlpKwEiF1UmSxERRk
29/Km/kR4lKstj3CzBTaz2DSLD66vdVCkBiVxfOww6+AQReNsVObMsLZ1zE4Ig28vINRmox2zmfV
/P8oAgaPtFLdaaBq2hiKRH3B708yhvt2Nkens+E2U3XM+dTzcV/Wy61KNS4uGJuQwYgX/jqWv3dl
tEwWJUNMIiKOEq4JAKV8YDOIcqTgXs6ZGTg/e/yEGdC8aR6+MvHerky5YrqaJcA279U7/jzuhPhB
B/JVmuOtDNyOnTRLecyOqRSFrPgqg2V91fDBPWIIqCf65kJB9Nh6YEq2kk/u9QNqH9LXUuMwkvPu
wI9CBFnnuqGWF/JqPzOg7skQSzfdxdK34ZySqzakAWq0Qll6j0cd3U+okWC+WYo7Y5+vNM8q3B+6
imIxjuuhaOGXphpNGlDDCkW/WyZCDL4LeKz1o5ew9E7bPHllwx89eGs5awV3DzQrGo8eL/lnwtdL
BGFLrReyVYwQeRA4uHf38tpQat7PqNRvKL9JoG0LdjwTWEdL4vGEnf9GzWOL/Fnb59Hl8MScxY4e
ZMrk8db9pJU9ZwjqJlGJOn+cNOxEWHu073ubNoqIqzIFVRnjHUzlz0qrND6pu0+b64NhDwcXgPVs
448O5/wL5ffUGVONrVYRb/zsTFNsZr7p7y+juR/xz20GlMbGrZvMnb39uoNw32jgfhsHo8J8IH6c
/jNCllBVqdpnHzEVPlC8Oh2mg9BkfAWbmueawcLDj/gkP8v3rdFjP9WuTWOOmiE6dVslpaQ1ar68
wfTJ3z9FAD1uu8ur4V8yFQV9AQ11FX9KNHrFeFXZib6jbfkaphRTDtKOWX793LSfSaQqMJ8UJSeM
BaTHjno95NBpeQV6aDaLlGdhwSr9/eGvfEfwUz75U1gH+RuYeIQQLPI+aNIe9WOLXInsAb+ebcaa
kDmsWTKnYu3k6s533mguT7QkaELz3lwHfCra7NbefWgt+WIu+JTAV4Qz3OpICP0G33NZ/XXfaXRg
FYodFt6x8yNXMyFWGr/w6uyA654sSVd+31OVgalFQxT3tKZ0+tCTfIaIbLzUD2t1E80pwZx7UJdp
aLcf+zJ2VUkmwdjiiSA4I/xsfrjbcQmS63XKKTgi7G20Cbpos+c89SKNvRe/b/axRDGmaCzMa/mV
nD0/3aLZ1AV+/bKj6Zkr2JJyDmji5wEDppyY8T4T0ulFc8sGFq3wENJEw1F+wf8gXGkFVt/OfU2V
0SJd8WeJgm+V80AR99Q+73euPuKbAKX9vkRqmR8iU65IKaG71Y2EU9L1oLLt6YwqK0jBFEqGPFOO
5Zo8MZI4PpLYCNSGlUaO3ALNuFz82INRKNslYbDzquj/L20h11qfiX1Ca8qJ1opXQxhNobMqqGRU
BBJt2umQqkXaPVScE8dx4IapzWPTeB2sXIorQzqxYTaoGjD1u+xdJyDCoe0mDQRn2xCszeuO0JoG
NCEvanWz3XiQ+a/lLFkVS12h/EZUh3N3sST3cnPo5lNH/e+iL2QaSHB/fVGh2j5anLryRiTUKSe7
RC8oaLGPMgmyR69RIBzl6Hk5i24uBDahwmsmmtGvAQQ+5vbGFAQ/fm0sHu2QuPythbimTmhYWMuF
oVnYfRraLpOqB3yLYar3SGvuVXPbBCtfYo/qxGpGyISauXWpUOc9H1tIVdVsJKtjBiazgT2YyW2I
F1FOpKvcRBEnku2TGxKpoqZ+iHkZMQeqdqJAqEIfZqqTgxsKWDMLXToGq42CWNEURTnV+8fytflX
i6HkB6YUdeG9zsxjMpsGqG680Foc4xUX0ZuBV0Os5M1dsziC/Lxq7zYAdVjEeaBLiANoZi2j94Bv
nU2qcl1U6ZvQ3r89kTlZjRC5Hn3wo2UCOTkj8X4NAxpbE7X/KNZfnw/wE1NpurrVHp8TeHz4O08w
GNcbm4r0ay4kT/aFOK/cbq8l95uaMarOBbNrrSBRv6y+URZL4Wc3vzKBF4MQ1uummgPFy6oC2S2O
o67dR1xjWGArqbkMvNgwpGE6mJpVmpeThDwZTstGvVldSGhkVuLfbc+ikNFXt5f5ZJjYUuhfmABw
bJGsgHMTOMpT+HI1+vCTpT9Xc/niLKEts5zqDpc5fzCXL0JhTN+zJRiaWazlUPPBXfvpcmKOVv/J
p9+V3h6VgIrWHbnEbhuGs1iklIlCwEDC2u0OtOfe3CQETxjth0sJuF39hKW7Ax+pZEu2TmsNq3sM
oigsj80hcdsCd2QrEYPLn7uFxmnhE8QenQ780RsOWk34ghVX5Rdvx2tUKeX3eRm43/vJSQPYha4z
I+0+7m6Xbxp7rCg/6u7kgH8qCQdBQMPW0kX4BethoT4IkdSg9Sq0+gP8crUVHmk31lN42WLHZXdD
YBAOPxw2A9W9+kE0/wlH/InpIHlWPfWnbJR72fwH1V0O6YYbfx4jCuwNu0rkCfTJzy3XkmbWucfG
lWgPOtjd0uidLVI+vu18ZEZhlohB78fSOtTy69fYg4/FUdnFKUyHd5TmjCYOSUCdozDonahOFA1F
MCUqeCqWykHUTC/8vE1ZrxsIPzkozhWO56qsO2M5eegxKMd++FKcTHwofX3KwqA1BwA1Tmr4rZYc
YWc7tEKE9t8G4OTYS4/ikVeoYmS5xXoz2OScO2EcFgIqeQd/B01egpLROGLQxZyizHgI/up4laBO
uKhgBK/bURzuBLMMHZfRetbWqOSGvNOS/wV2/RjYyEbofCadT6qE6/PC+/M1l679dUhWLsxa4rb8
nX20/e3UnhuL3MCPzg5aw/S4QqBcBI/31ZL8YGJsyS36ilTazAeB+tH40oHPzd3+7CUMGxou2at5
4T0FB4/qKREgOwe13rLBO+mPCMOu4OtSBZJodWaqLO2m4WGYg8WYojBGflRQL7uTR2fsWEYzATvP
RdLpgbQshcxTp+2DoluzWuVyCmPaslW8D3kJpGk+vcL2GF/MhsLF0SJICy3wOmKjCJKlkWybm+oh
JQmlAfUNUNco2oTWNadLnDduSDZjpgaP4OWiFL7NJqdUyQpY47jhrkkedWun7BPe/FuANfxkcxFg
ENEkAUZLA8auo3qXZzrYXnRgdpe3ZKstiK96MIdMUnNvldQvsywcC7XjCyZVfGsD2+lTG1E1ObD1
1eD5jSGS19RwGnPsv1j8eAsu0zIu/OjM5AQ1dZCp8JNwXGAa54tQkSWjFfwTRi0mKWPZuesgB3/9
QJHyujmbzPc9jf3nWsMXhYSyygs/IATgUz9idpKjQDpEwRBCe5AfvNjhCdBKa+g1FJtR8OPg2Hob
lyqhNvxsUA04bxH4hYAiqn4alr7iFbbiOgiiZ7KZMMS4kH/03ptjdeIDmT4Zf/3fZC9zdWM8xPZk
Esc0yQ31B79tInnist4sdwO4rFfZvK1v4iagQ08gjZ32zUpoceiavAe2gzjghXG4G8+nH6bTFQCC
MbN5Ax2H3cS9Yt2+HIs7O04SVRLx9XkHCM0i5vlzby3hH1xeAWKh3i9Vk/x3SJlZksnGQ/dBUP5j
cGwTKL4eKUeipX09H5e5vaIcc+qDI4bShVDMuYovpT7gWAv7OxTmoKVQBBpldQPUsHTEVgEAUvGh
avkI64Y7ab8i6icdGKQHUVEdSbVIEE5EQhM5WSauW3KlqNtITxH0TXkdEO6BKSMko7wb5Yp1sgGx
SrSIKnrcYKHorMeIByn2HOvjFxQQNKePbtJpaZFIMTb5dbyO5lN7xDb6Hb+F4nx3GeU2hhyDGO6y
+yNGCQI3OHoJ0qMPQyYxuS3gSMGWHpeK3irO3wQSe2TeqJjVAl0oHERppU4Jy6AaAXvtXYifSR61
V39LKJqO6lFSLwiNIWPb1UMAlyWbJDOOXBWG+0bZT/b98fxrW+EeON1Lm/VcxiA38uo//0+wPcJ/
cWDm3cdPk/eYCrVCrUeYQoLEPTo53WY5wr9Vc/e9sFRGBPziFAJmwdOxuj4KpGVuXL0MGOKsQWvl
hFQ6YcpZ6hLJh7soSU4rrZgxtNO8Z9GDZ7mnPhGxFIY51FPYJR4Q8ppLHVcZJLvE/IgnLKfQls6D
1be1i+0bQeMjC3xllzHcd6tvZ3sv77EJJruFyNaV42hrQJ6/8w2bG8yY6b2l94XhB8gL9WxcYlRX
fCYLmLa+0B+e6XkpYVTazew7jP+Rs2sXsPkU/IUp9c7nVLyyneomaRw0EfqwIkjyaDuYvtBGEMEH
X90K3FspBpgnqcmx3jc2PbD0nDog8aDEPKPkxxZGYzFxD5nrJGwvRBqxYHkpLPFurDdb6n436jUR
Rv+veHM4CuKkQBGl5spDvz0S4gnqKEFfgArjb+XM0ZI3MOvHls50gQ2alqe7oOZpdXXZI99CM8iC
yHi2FXOeuXdIVOz0SS/3iJY7oXF3m29sZfeoAZFX2l+Cn4CwWc7wNu77sR1GBpR5So5Pj2UoO+S/
Rwws5svTxeX3k77XtHbnlG8MAt4pF97kn88sjSE4V2P83pD0jsNJ17CuTXj0ru726jXy3g+uuUJN
d7n6WjrDiB7rBJZBX3HIKuPmI4sSoJi7x2Zj452JTEJzmuaWUe8ZZtKh4GttwzAuVJysxH2ansAr
fn9FLfd60H9UWBvPLMQ6Md3kGNBQEeWWqf5rBEAB6wDnWD8D0jYN6lCtxTdRlEVztVZkLdK3e0yQ
DZ/D43rIgwlVoby0Hf+0+dApHxe0Xxzdw1nOT4pv2EZvYcsPdiehcFP+xXhy1kbL9AbSmczXlqok
ONTaPXFiWJ1vCqbG2JTw/2VEy+EW10BPnSsRAaCZyXVvsyXfldUukBa66vV/2MxQl/9oagYoUrN1
VMygCThF57+kJ+9jjf0bIga464hafxSwxJ4Z/dkSdhdIb73l03p+Bg+9CWGdyylqpotvdWrbSlZJ
lck26neoygAQd0t0h9v0fXnn6AkS+nv9ATMLJH0lnCDItz8bm53ofPojKK6MxPsFbiRwtf/mdhTV
oqPXRMSucgPHq99MTOQSEWFIMg07XGMeckn46cCvcQa2hNxC7AF4Gqy/RDysOjaFlPUChQ7rZ7cj
q3PQI5+qcMCFm9UriJ8tSps36GA7BZWjDyuZ04Jiz5yJdaEOuJKDkDdcawZm6FnSf/oNqcigGHxz
2kRE/Z0nK4QNsXpySm6Jh5hozB880GDeNzJKfXhWWr8ckWT0stjtUHXRJSahqGYIdtKNU94HxOcS
FPd03InpyCkOEB+RrfC/4dhWoITMkIy1UmgPpbNYZfjqvPwO9leeU2U7u6gvOvMGE+2RdvHS9P+t
thRbbzUZAUtu8E83Zs0qQpAGEMA2RFeOkQV30z4E1IMjy4u8A6hFNS06K1t6LmGXNzJVvJqqHOr5
VvpVKfja/xYZ7u1O0pczZaM3Om7wiMVUdv7+5iq37ezYiWqABh1JjUSaVZGc1WjlyL6JuAWsD1W4
Mf0hUXEPgpQRI2WZMPrdFh7xGnvpdoqbmfJEt2S24PX1wupXdrc0471q53uaJ8be7djP6mxCpLIP
QGLIMJzUgCSk4NRPfeGgbLvp/EN4ijtikxwOZNxmvDAbbnoLWmMcevHIBjZqPMx6dOgm9MYlILxj
SAbiro32YGD14jQzELKrqitphAbAC03Y3MQysIrJTHpLCxta8dRmB9qSfAwyT8Oi+B5s/0tvPPgO
H9MKLIZWKErjVAIg13otj0tIpricz125M1R1VG7osVZFnXytGlIV5U0v3ui/PbWywHewn4eenEdn
7qFoFcB6yZCm1PXZlmCZL8biGOIHQ8fNa+KytDXdopaMQgWsE6rUkruH7Sksb799aPLIWqAe/4Iv
+r2dFsmRy9F8t5HBhrlrtsg6SBOXABOoVEiRfGvWWYVzJPnrqtdDb5Y5dGwVYGOkVDj1H4BNn3wJ
ZNpea1FY1FtyUEN3pOGQAVDnL25a7hpJlh31eNKTNKGQL5E16/24INfrnYR/7pit1aZmnJDkaZb7
fHmsnAWXkqm65LV71VDBAvO9vQtJuPh7ntPBdFj6Dytkgo2hLAxjDO1V1npeWH7xQYM99TreYoeO
E/G9JG1jd/BluTstEO4RlWew3s0j51LfPjSgFCWD/X/tmQI25APuZv5L8NPkRK5r8dglUvKYvNHk
jXQcFxXHQdp1aHJSjB6SThjJdKY8ULm072r2XMdNyiQqUejCqZYnkh9OcuNAgoes0sskTwYjSxra
61t3T0tkvZAecrbMsYhi2FsUyhqM+zkmV8D1/aWAjUFm5/llj5LZK0xeZFbThO1nhQXtkiObTjZc
epOjKiA5N9QOymnDgh4zeoI4KQq/I03Wo3ae6n9vttoJSNtHXMQ5mvUm4Jij7cUa82wapTppHHOq
AiA2bPrpysqEtL3SIU4yznoSlS9eNa/g2K/V75cbwp/UAqcMIHpD/brZyfTsJ1VFEdDBkTr86a20
lxx0J+/okm9UO2XwXjc3q+wyhN1wchucKlT3sz6mVrw1HxawA2N2HZYjj7qt1LM78kUtRg+6iYhV
wTWYdqpTMz8VozzIDz0C6e7sNMlsdhWpK9NXrE0UvkGANDAg6hTddLQGye3QwTy0kK/JuQfrFM2U
y3MKPXSX7/3dHasWE8cS6aHU9uOoE0nNKoVuCDxxg7sYjsK4rquhFruLf+5ETLwpgabovtocBPtJ
YCPoC/RPf4IVvLD6R6d99xFrhHXImp3PrVliWVNIqEE74UO9wwzZZTS8S37sC6D4JqZlwLrLg9c0
G9NRmksyqkS8wsrKaYlcwKLF77Bw9MZL1Emz47NP0BvncNDuyNf0Kk+COhGgzp77og1HSH+bz2Hy
7/wwDlFl2U+B0ZbisldG72riZwfp78mbr3rnchmVwDaNTitMdDEP54rWG7EYnNKd7bKvqlZho3CZ
dPYl9peYZgQSpwglyynC5+kUbrb7tWNJbSQFi3f4Ii+c+baZyDO+ocuqKHKLpJMPpXgiLRJlNqdj
ZQxFBXE4+C3Zj2Xc9cmIqvjYSu03MBsRb1siBDjhHzZgH6FOV0mmiRW0bbaVQzTnPylZGVdO9e2k
RNKuQYSh/zs4u292y36sWGkYd1h+eZ9R8pKdBu7P3D8HWMozurcpWn6iI3TWIhL+/p/SpuxkNi1l
xYTZ6hmLBx7ZNd1Yr45Bfr/RP6f7bLzJnpc/zm821GwGn1a/1MtsBcLLjg69Q0qEPybRZ1k9S/jH
eO+L4/1alLZG5gED0Dm6ZQL+kzByTg5Om4QiO8EElte8DJudATX9EiciC0KG2PpPvhDnLgSa1gSN
RAC7UWoTKjxBVzG4j1H/Iut2AoG7pPBClhU4aXPhNDUEkJxKXfnfMN0aRmqH+HcHZaMWd6aoSEJ4
LnLixw6VZfLsud1Kv8vJKTbN6VGES3PpWmZGdfhCYozw1l6KMoYdf0xi56/85Mm2RwUCoX0CB35p
xN/xML8Buo70O+696lQdIGahObJ78cLlzBZ0H3YlAxjS1I1fS5KfjnoK4scwXz2wUPjtSGkY41K/
tRMzy3ugPa1haRHlRjG85oktxK6nhuzSttsS9Ie+oF0tl/7z+cyjRU+qX3S0ondjvP9E0QU9p37R
BJOFneCNLCNkRgTwb00sPVOqml9vjdWC7+XvtyUxdai/HDogzEatsLSiGQPJCqdVh52ccewm8DbV
7tZVyVtbNvALT7c1q+LihVgxjh3GD2mEJD1CPErTGWLs9KTcBSJ+as+XOL0PWtJ0kAKNR2/bZ8W5
Xs3NbXlHTIrpqrHpvaqT4qnJ2R/6uipIL6oomqy2zefI3qk+Y7alartbiDNq0W6XuCc697Qe3hKD
jn5aw4WfJondAIbeb/YOTEe+Hl9p9bUBnRm10r9niXqgRYv2VDmaxMbBNC+mM1m9hWctxRg/WrGO
5x9y/t0T9WBE2QohVlW1fdwD3KO++ssQub6N1mOjpPKUH4zkc998d48O2KylCvoC8oef1D2QXpCM
cDsfZIeCmD/oqwCehr43qF0qKPUjwwkHrpU2A24a/gxXV542/yCl7jVrY52FsXwl1cpARGNkMonC
LpZ4A/xr+o0wsE8CR8MDgLDOhHRnZ42ZFv4XX39ySU5y4LszA0shLmOvW9wi+eR3jivgfjhd5ukE
WN5p0M/7Q7lrWPjOAPA75tfgGmUCaFbcPZNABL+sE8k6wDyJCYFhVkguphWyrS5v5EqsqTCs761I
SVDutEj/IoES2oQ34uswEkf25qH7LnEMuUPiA3J0W83xDaKImh+jr8SKS4y4FEQpf/YTLUohrP2p
CbIKImQpPMqdmt/8uyEFwyY6it7xxjr1fYK+6P/OsBTCuFbe1aBFgNjJA09+i5dfIL56xIrgDFlf
2Xtew5L5t4GZCMwVA/q3bbi24QdOkxAQdYq8n2ATKgxoD/4n2qqh0VAQcyXsEoro/jPRjHdtQlOG
wusWD5cZzVSJIl0jLPt38MXBeorKoAcjw0XLlGtklewlVCwS9ts/nxZvP4trhShGxKm06ktuDVa4
OreF42Da7VEpjghXxAm0l7ueVWviq1kyVtL75YH/jo9MwLtLmi7O7VZKzeOXZjVsASyg3wTwlKma
SQtFzrmSngHy6MN08kd612O8O5lju6e4uSdTNoYWa8y5JVzFh5Tv65svgzXr4zdACALhO3ayzbyB
z3EwmtY7U5BRGHd+aOkBiMTipdz43PyU3XWGxcv4H4E+021CmzBFsHj1pqAnstz3WJ1wOaKIUyHl
jM8oqom/GecZ7d1q7Q5NjssiWm71vx/H+XbgDv21HPP75+LZpQ0hOchahOdb7w2X2oPvgfrDj34G
2TRHIs8sKtrZIgXuQmOcCQVGGYmHC5KW33cqD/P7/XNVnnmuAL/UMyfdBT7Nyw7QdQUzcKepzojG
H7YXQKt929HLGDaF9ewHQ24X5UaXR/ezZulFlTDMCp1yQqN37AZLIqVqGFGXJsnDn4xCkKwcddrw
AjJf63PKCN1StN3G9ksIwrHLLaPGnv8o9Mpjy04r6nq3KQcreB9B0HKPZupLaR+5A65NQtRz7bOs
tM6Hl8x4c1WS/bxNDOjbmnqfYL4pTqR1thCwGW8IO4HCYVN5sJ5SgMLmcjvCLrCLLfLtLLLoUqU1
OazpB+rXQIvKAaFbN2Sa3kh8Ysl6hQ0mu4biJXqlzPCMdC5xlZ6Ilb9uaLrmtWnKbE406ebLZDrv
FIRXaIpYR7kK4BqK5wz6+7OGeftd8s/sHI5zl+Wlg8yu+sE54N2K4dPMY71Q0lAfpUz3FdWHYtxf
we68eKwhmrDoAwNVVWdx93zvil12/GFVSU3DZGfXwQMxtsQm3GODjyizPi/BdRNDOZcMuLHtBkQy
Z3LdW40vOdzTXKjIU9GZkedpf2A0lRMGbcgXM9AY0YnafLv3S2i4+kS4BRgrjPgfhmR9EL5QBvdb
gEkWSCC3GfhMgNu+2yl9bbBxnLllBRXp7FEmv/Wpokfzy4dtiwcrgRd8MULdzfHWnHgXqakiOIuR
bQQzkTinQelO06iNTFiiyGKbM4rmER0pMQ942Tc14e2mIMcD7UkslMZbT8C2vcBVmLIYHnU487LI
OUbP0IbhO+nETkID+LLywxwZ13xCxcuuisBUY/7mnLoQOmJhBNSY/eAtK1/AtbzLxdd6iz7Nqkhw
FZvmLHCLlknycR3/Rc/30t/HtxTj3VgeviMypl6Pf9WMl6/kypFc7zg2B5tFJsaB1JWz1FAfOWQB
Fn1T/lGRUhO38NT5tcpz3oKoA2nnwYHyP053gZTdFDN1IgL8kbljz4TPW2pHtryqjCdei0vEzKUB
kuD7MdlYJ0ymrruZsDNT5mnb9s6SnGHjowAaxlmyTsrVEwQNBOmVH7oK0vTImTOBp7XVyr6K/DYy
i0xMgyXk1niUWCiIZxgM639PCMFKvfU+nex0JmuTAE/5v/pOWtyU1ZNS6Cj1yOq6aWSISE2ly+la
t3HtG2UBv7IkUqxHcBjRXsXcC6D3MQ64wpCOXKz9j2xmG/fck0WVaPvgWWXYbbICq6C7prAWKYyU
ZBMpr2J2O5aoEcqgAXzQi8fyMz62p9cr22blhKIpBRpLZWGaOheIFOW9gK8ljmqfdU+S+IHoJQ2g
WpYYrIafCKIOvFvHaJSnHTuZ50u5yYh/Ful2x71sy8FjvwiqwN8sI9twZH/HuydEp44ZWFvSlJcp
nrROjFg/Egm7d2jxRL1Nw5W0c1CM9gS/2f23bCFHo3Pm6zeNlCLg3OIWON6+oe5wGkXf+5OIg6Wb
DJnXbWATszlr4XRJ8Tu+TQTYWVauDve98oYTNYDHTVRnTvYj+AXxGyVV0LzGi45x2ox5jOzal9Aj
hzz9ThCtn1LNArjm+6jwn0vmvfGW+UX1S2W/HyHhvmD4/uVDYx4iCPwyQOxwidf/vv2qsSQnZMXu
koW1GbTXvJfRfCjojrRBKANHn/kqy2DhTFjZQV5rK54HCeVtibvFRJY4LJhqCWiivGn36fPeNWCp
njqUl2XwpnADUzJh5FhvRbauE/mAbv/Q83lyuZpoqbR33ZOTI+ubuCSXoOYcrLRSqCrVZGCD0tGt
CPHZoJhf+u9/gOJehRYECcI5VKczfSOBA9hCm4SzuyR0t9qabH73Irh1zD0+qH20JqtH+tpoYNdZ
/0U5Ms4gFphNtb4NymrLLMi3OhIr31MlJGmTGI+MMkvvejwqxeMa007/5XUCaoNBmi8y8eu3dKUE
7wADnYZumpFPG7LvB3akWrgl82KsxGTcvA9bMLGe6e68sLBA0NdxKEaXNJL8xBRvVRE+/M5D73KP
YsVE9EvWepqowExzN4p2MNZUeNXv7hDV+eimvmJQdiiXiyJjLnrKH30f9Sp9QaC7h2ufhBUEutZi
arTJNwrgV2Etv6ceiWSoZj3LB2NEMbJdOTpMzex085VeCurRVyOTxRmnFx5magSrc1oxBHbSUUy4
fPxD77eyGco1w88yOC3RpgVmgC+FqBRi82n00GJ/L1/rQC37mFdW141iAmELphiICxHpAfLXXFA5
PJ/loN+qE/quKWmKbXY9ausjHFyBmTCddsFyCCo9dd9877o/UC/Phq1sVaJamy1GWKQ7W4vAxw/9
/3pO2GMV88k7cv1RJ4uPZQw0wX5eSdpLO2SS2MVc45uN8FToknrmpWfYteV+E25D/7iCqLwF5LES
uGCR08+MAM3s2ppLXi3W+TiLMwJ1lq8L7Mf+Tq5T9ismHapj9d023xjk0RPzCupEosPulURR0dMq
6hn9x9q8urJt9JilTHK2UN1SrpLKlId/cC6cQKvn4vcxlUDuB+w8nlsAAg8NeFiZ6h22IIhNtTw6
8nX45pIFZkA0gLEd1iDcVtcGHdSMJco4UaRodbsPO0SSyw6sp1sc5Kn3Jd2gnyuQjml+PGZmlCsN
SINnvPnIhfxWulb/euOevdtO6GgZ6kmV/5vmb4eDCI4hg9EfA4M8GtBDdLKnOwDXQzhxDCVVj6Xw
LzQ/NoywMEal3EL7TtWjhYk3JTrgTHyGiRcDEWp/HvXXwK/Qw7xJMCgpl6FFYKmVV8mbd6hEhBYk
7S+VvE/tzi483J+20AYA5nj0P7cmgEMWiNvfkgKRi/YOrnIFl1NNNDuBrNEz8MtE/eTrbs5riN0C
hESt/2IAhF2aauY8fxh/nDWjDZb0LeiAUMEuty2kFH2ktv8MgWcpL2vrO0EacedVmmoFzBLBXYuf
KEJDGKavUpG74BN8C4OM5ZpIvpEBSojgTdRuHotBBVReavlzF1cF12huK4Etw0TsmOZwuhh/cjdj
I6ZRdXCOCnDwQtU4jYioDQfTQR+P7uDtqxddspBG0JxuHPc7oPJk1O5vYi5Mp1hV/zIow1HdhBCk
OBqlKGzEAY0GcVLd1t7pgRPa0DqOf7UuxoVGzpb0pUEJsapBQYH0GjWzPcd4AWZmNj5IYdKLVJp1
G/Xy662bZ9PGVm8AXQ6U8Um18JT7ZiKQR8geBFPurGByZu63L3gqv70V5579FFUOnDbMWdNpsBLj
q4Oxq6atHR1GIzSFT6kMAZIkEcNSMwr0fyiY93uG6NbSs/dKanYtC7qOMHe0bA+uLFmG2yf9SkdJ
k+blSGGqANn41W8v3s4aEC1C6nilM6MjVBjp+smDOKtyp5kML4vXLbAe0D++Tmg3eKJGjQS8e/Xu
hn0OeEDTY7sRgWul/+0C3gOt20SFj9OEKTw91WqH8EzsFQ7TqcvA9ldwLYp+LzXiV8VvpmLg4nOa
E5FLCrg170pASJr8Jcbtt1GvUXY5UsvnmztloxbJVtmb3TvW1XXd9K7UQoZYD+NzVw7yhjJAElj8
SngsKWW0+5405auiQtHAAAXJy2xjwRj1kxAbNd7wBiGm9OvA6w+2dJo+FIzIbFwhEWtg2QUUJKBW
ykNGnYHwoLtNDdp6/GVojs+S3Inyte6tqjrfw5MtZBOwXsO4n1W5o+wdzNrq9YY0j5QIKvgVo/Uo
0FQRZqtS9yvCkDw9OYDsI2B4GnDlr0Hl91ab4Ilgg5mggwVXetqZgCBLM0/nhKvcY81v+pouVI3V
bE8iiXaTp46Sjbm78/Gm4MCqI43YLnpbx3uUVPXBfBNQ0bL12shy1FXE1rpZ/6r4DuIWdQjyxLc4
VPMDWO0y2efMDZwhgS3mMo4SNi6jufPpZj7NFASWBcjjnscPvW+gQsj13pds6ZztXcvFgpbrsErV
sqDv09bypFdEjTna90ViEhBQRIhUSdurQaWSxn/vRYIZWlia4Ti9TtI9ebO+cZ5L/KRjpcO3SbUL
B47ULtTX9L2PQOISLK4XOJ8lc+51QQXiX0LI6U/3hdMZhlWXuP83NclDuwlX5/q0EiOLiU52bRg3
OQl0HJknYJpO8hatT0J7YXqC9oUhqPotQESOgjXEz53H19FO2JvUUguer0BniEDd/na0fjFC0S9a
sVz5uyaWawJ6PT+hv6+ThnaC03cXV819Bn6JM3eqdy+t9bpGeyV7S3oFVLSk1JQEV+5M95YBKuNg
uUxSQ71dW1DF5Wh8z3+HA0m94uvsWxvucbgw7NsNKrR2+3xUTRaxpj4aMndNCtSrNsi4gmAQSjw7
oGo2TB/vT9WzQA/DcjMeA/LKpJbYiIH+pvAcae2uXsgNV1CM0EQSXG8beWXFpQXBEUh00YaWYbD0
y++7Nj8ZdKK4JXPRI3xWzTFvEKG1BHuaEuCuyD67v5VdV9GVhzDuHubt55hDcNbdQPrpdX00wJHt
DS5xSe9lcwYwz5drEOPyw1ibJQVVfcX7XSVATzanw592/qtievseJWN5m4DrTm6Ile48kMun8VAq
bH1+iDOwgTU9GW+RdiQsPfCrYLR+eqrgbnhMyTq1jYrbCvlvC7tlV+B6EfiUqoMQoTa7zINeNDoz
84EGbq2GJs7KzEjV15fIgaARkjLTktJ/vWYoEC2xV56FJ2ckXNAqiO88+EvwdASLa1yh/y2FUaxj
SF9dmPw0OkNcWGcnoUk2x8KWvnEhxQYmeyKfGHXLyfBt7e4Xnoq/qIxrDlBgQMcqtlrTU2XY8wGu
A6etdzMisgc8jK+RlIOV2yQOO/dmXw61KP+SDNSfhPlq63na1iKP/ZuwmKzJ8tZQOaebR78ftiz/
DX/lR9cXv8DNbcrCcyX98jeluSonpolBS3Xv8PM4FbeLzMXCO0N/EKHjhdAm40NIQ0IkLUSIxbqC
PCD7bLibdW+AGtEkNZqPj1FDVF4x4mRi+aKCkw5MoTQ7tIuSSPMOHtwWV0L85UeR9cXaay+hTLaN
kGj4LCOeGqe9+pXYzp6LgyhquavzjchpJGEzfx0fA9PtBtUlDS4PmzB+kFUS52qZu4vVpezXaarF
buK593pAo6e4EMeyAmsoZ2fL1/0LqrfN4WgvthHYD1Oa82BAFEB9+yYwjE5iZz/U8Ve/oHvRM3Zm
7/rTgurJMyq9yYo6hsdbquqNslk2FKxXN5+5MdQr1tg7lrtwqWQjhlZGHQU85NBUShHVpTiCEytv
nAK4X4VQHvAwUSRJIpX1uNlm9l2N3UksukMXsGSb01pCVtC1BdUL7MwJKhVLdn+6h9UeXycDVVuZ
uvAVQnOG3rgwjO0oqcKEHA53Lizf86SfOv3jPKe5VXrMs1R3E4BTxZhaovmy2lkefR3k4b7sFbqo
AIT6EyiWSy4ugIWrUDow1IG0ks/NbVrkhJ37nVcTE4QEug/j4oYTWnbhkayxBhss9eJ9SvzDWqiA
XyT/GihcAqWNtLYJSl6CUyUcOli8laP6Ak+wa8UfEW1mOnlcaS61fg9fyPb4BiddTLM8NNop/0Cj
5cgCGG5NhA9KLofjFctnawaqTA/c60FMUiVuGdyihW6DMFGSr1caWb88JIgKQinOkGh+ZXmsboG/
Y+re5PWAMRHTfba0U4DBZRLXTAXbIvzFqR/HqMwBW6v4LGmU9X/81dx8+X46+MvH6PnEeoFWOYn+
s7y5yS6E1xPKIrTB/TmVv1Z0iND/NYgY37Z5wNzF4PWieqwlZ7h3CPtlTySxlJq7acK7SGB0bsDk
AwmJapUsnV/n7nUeKDw8ZWLVsi78jXbmpumPQ63Ge1B98Zxr/22xu8Xj4fc14s1EsISTPR7BNHcY
G9TGyHYtmzUhZ8BYj9Clbj/wc+hsDurIkOeY/4facH9IT3OvoGNlnXMjkcnzlkr53EN7Uwm33EJ/
aSJAEU8SOxi3Ej78qcgXWYwbHVe0VaEJzs7rlGEfHiIhp6oSZREJb+eI5PSRhcFe98N0YbefC7u7
J08qxFPy3tESvJH4rB8l047KzW9tLEkzeNEKJB0plYFS5C6uSBvD6NoQWPgGXRlUy6FGhJHZYxY3
fV97eHLjbwY4c/o25NshC3w1phDGPyewFY3/nproz21GhsXPyzcsLY2oaWyB7z/4BQ5FUQNN94ah
PD2vvWE5xHrsyg7OPnw94kDplJb7yjrjYsD4ql8aUCocpE62IDnhMI7CX+vUqx8gFccNo7p5KLg3
zNYX6oQW79mSJMgYXkAnBFr+jDSUpCrG+FqElGRPYwkntf4NmRe2n/sPh4R4SIsS7JCQ3U0nv3ui
xtO5+gOe18leyC6866d0kWMEsuGvJPd1cp7LVZbudK0QDrObUu/mwA/IQQB2uMpRLVOk+FDGMmTi
8fzvlBhTLyX6nLKR5XFyJfhRcfpCNyUR9RvEbG1RXiZ/ILeTIGJvnTmF0sbKYSLkvcwa4L5Ex+9D
N21epJ6dQkxcidXrvz9j0fEPOXwqWGmgfQnaKh9dXZh27tZ8+YLWezAmQkhgPOCdVz79yKfFzoTi
A9nSgoCeprutqVH2ybS4mGL5hR890sk8D2giH4gT1sBwoJofursvPRvPNwMzjZ80EJ8X1HeRzU94
74JjVTXrNHLjQTv5yyMuK3WwYJ3Rii+SeK9LeSLHBJ25its94fNz7iqlCFe0Ga47DI5KnbcK9E1f
LLMkoY6hI/52zU3Wwbx0NJFX1waqkS0CRlKcFjqcIY0IuxJnzdfpIEDrdWym07tFO3AvA2O7piea
I77ZYYUnwLUW+n5Wc+ArnixMeXx5/nhDfV6kf81U3Xq8cnXSZ2O73JkKQItkgcAYRqilIseVtQJ3
9ViFQw2NL9jGGWZadeIOTD+68ATci3kaow1jdXYKhc69zmkTWiVWkQ7TvihXAZLOooB4Crxe1sX+
62egFmE7YAwnqzM5MRJiAg/6saZHvqz+XFmLa7Dr3j2NNvdLpC3YLFpZgR1Q0KLmQLrWeQrQblBr
ApaF0FSjWHytVr5Hi75gMYOC2j9/zHuGD2Dg1W3SebCE2qiRYTZbQKi8umY/uUk4dU1DGT3XgSdW
su9k9+yLDGJUySj1UDCKcj2K+/kvS1eqKDek3eF+cViOqY0ZRWz44/tAhN2CqjQSvWzCfSGgkkyg
mPOwJeMi2/bAfrWXC1thVQnJ2MX7clBEZ9pr8T4UtKCVIcr1OSSViZmcrG6SmsQ3+i/smUxtL+4M
jhx22i0yJX/zUmEPh1VD77xA2I+xkRJ/sWM5vtgDyy2tOcV6iOeyuoOqMEI/UeKxE9hBHuP38KfC
HxXGyiBbWrQfWoYvelrtTpTNlrMtzsohNd8YoSiakRU2qhpckMMEqyiIqdk2MFm6oiBu9W4u7KuP
JodCO0bZnaRs/Q/rFU1d4KzXlk8uJ8UhxnN0hSuVpOPVYkl60tDyo3Y72fSd073up0Xw7XrRrrqk
s78V65qe4P2hAwp2EzpNxI7QDVK9PylLHPavLYZYVoHGxzZ1E3m91z3YnNjLAse/Zc5U+Shwf8yl
sgpAIJqk1lzNsLEIyUAEHsI5TISS01txblSFcvjjVgDj8YRMMyVmPsaI3KxVHKBPFyWPE/dNYBuf
GTpes2+7gjQ1T/DjCXi0cQvjMx+B6j6p6eqSPaGYStaTSVyNixGFUAgqTfDcNjqxQw0iOWt0/GYG
dWbX6gxQLDVuuzEWAh6X1LZCftzyccUrG6N4wAfg2Z+rWNNcqqeRHXfFBobdcf2Gc6PkoliZWzJT
q5ZZesbeJ7/n3aZOBmh1O5O/rC6guH0a0eu60ynuqb9az//xMZ5W1aAnvqUw6JZHQ77q0F007PGj
F/tesv/JUBH4uUg3XAfRT1SCWuHdVDGwKlDGfdyTJGg4MkL6GLcdmVMDZijLoIOVsdn+Kdw6D/+B
8OTrFQnsdmza8V1c9zrpr8ljlEG6HrLWZ2VZ2LWtmzL8qLN/N21sFyURA9vD38OCp0VHJxPrhdpk
4w12v3+kCba8SUs9YmWpQ2T9YtEb9nMOTET9jYuJwM/1oV7jDKp9fjysbX039FX7iSIuYRt0OLWL
IGgWhLzjA91D1gxFAE+4EWjMxtReHit/8siXior+qgKfZENNz97Jq+oE6itFRf15eCV3UNQEK3sk
BB7/Htap2LpMcazKbBN/PCWHGZmbAJ+ytyOD3iaKPpF3MuH4Frro1jzLpEsVKdz9Na77a3jC4OvA
Pj4S1fdHxqKveaxsksduNq4VXrcKAgvcZ/2jOyc0XWr2HW4yl+xCPzz/Sy0c6XFSz/GRXbkUExZx
mIZNDbVePuN/PzvHlLB4HTG+DNENMxwhYRb/1aWcwDxebqxSdkvvSb4nNK/Gbe12PkneSWQi80bI
E72UR9A79wv6KAcj4E5T31jIwf1bq1zkPTo47QuVIY/zsEAb28192O8klbO+n4nCXSqzG7zBLRny
nmRwGOsjXwJZG2JqHqz4P8ekpKEGyWicv5EmaAR1nZSaLyZBPcHr4AXiqRbRV4epDWL/pbpwSM2l
hDsygTxPXCM4mzdNxQP7I1mC3n/NHeaK9t9No9i7h+Q+OXVp92FfDulFuINnvfQlL0OJ3HKpxySe
4hcvFVkNdzKRII00uQNW8C7I4H+XmoMrm6ZnyrcRb9u86ex0QmT1iQjEOMuC+rV2D4BkrKpXCkpe
Eo9TyBnEy1i0L/pQyJMHt28iLqMnS/gQOeUAERbmC9EPvCf22L1aKbQXcAeMV3QzLf3Ca3YQCPw0
8jNoYZf4twp7m1EP5Eng+Tu9UNQ75F7BzN1H14sfr2F+QV3q4YbQSE7ywer9U122TgmZJQs4jsUE
xjJBd+5s/hK1UdPH2440rXeA3q1f93WhVPB0INuPrGroxNDZoGBfq4hhNzWUbX+cU8qFAB7C0c6X
uluH+LCvxMUt5XmB2fmP4IHn48ox5hLcDm+g+0m9Lsw+DpLAgB6clcRVcoJaEnJYIXedJD6t6r3f
Oh0BcZf+ltC4g5kH8PK91RrA80/uRCw7qmkDnme3IWe02cwdqkPDhZzkoVVXugYqLvUEZgafG4aD
1EGbWa0No1HA8rW4JTayrClrR97pJRZnrUUQxr9m3dIreCpmwQxTGyPEkmoRK0FkH+YvKQ8fHQN5
3IhTPS523EslHe/IEyDfuZfRhi1T4O5//Rjlv6yg5n3P5mmF06KPbv2n8gW2IoGeFga3/U7ndv7M
+vyywnawIy/fUYlaB09GWTivp8kaKmxrheZFByn/pK2ZCgFNWVppaX6hOOacTzKsOg22jx3hcSgJ
vveskCe+rYIh4L0+C4PY3QXb/USZiMCuDlsVPwRGcr/77mMESy3AVz6H4eJY0B8uC/qIEgS/2/XR
sZUMUzx1VioJgfBxTGpGZbmCf9BvbF5kcTkB3VzlbEj6uJJdESYkewnk9Ft9QKKspvh6h1JTKLt2
fnEIegd04Zj6m1Y3IMOcr/1Op9TckDwfwALqSMDzQNXJfjOCxZj7FvShSrtvyV8df0n3ewIx+gUO
fWuSkG1HK+Qyy20nW3PfyO7yXJdu9UQyUNEzvOU1KK/3RlbhWssRduaICzvCrHKO/SYiDBva4g/k
V8qb0qIZibSu1aAmzNI2UtUupGPKr9qT6B3MR027+51l5Ps0NYFI2NrJeAqdDT8iggrhPr6gZudp
Fn6a/xAn5XsYUn7ZZKM9WdfO5w1uUNmkj/EH1cH0tH4hDJ/E+dyzYOG/V4N1dbPXBZ3xdOP7rJNo
TytURmx0RmNjJVB6xwLZADJ19Ww4qATGjXU31Fy6q90SxNYPt5LY2k6cqNponVDmbAlji00IxVlH
HTUlsTsvRvt/sNzEnUlwaKIW+PWB3iRqrCYWESm17yL54/VbHTfkiPCqP1ykpEuZ3plsc0nYVc4h
L4B/vDd7Prr8MvbqiqUmZF62kwCCfePkp9jqhIx6Z7uYMaaZH2et2reY8X7dzJ5up/fXviW6ojPL
Rec7spq/OQqYDRSWY5Y2plIRABtm1+VGChUQxhHrNi9yBu95uzseyelE0OF4Iy1FqPNqGFR+v4zh
yTGXi00MErJ2RxwZMvBiwEnm2wf6dxPajxIW9+7rb4IhPuOu+nuqGVv1MlY25+p0vzSvq9pn5wL1
8Qil75+gCXH4eg+uZDAtXkyYhsmC4SfuZIQDwRTRg5ws0LXqN8gWlq9MuWo4h0v3+u4GCHG1hxP1
vI7Mm2OmnXR7R4Q6umCHk1Xmjt2rrZy3RXzL2/9XOny+OidUOeEH66hGaxeqC72Zpmcu7CIOLHr0
0SvNc4ApA/tbwqIDsXPzQGWRXlW3y1JSSJDCBNUgjEZuNQbtry6XBWqpB7VhiE/0JOS/gEV6kMZJ
0VbUhznepN2LT/QnVwxgG30iDHm+6ZOAQu7P3ljDKTJRCLbmtozdgGi+ZG9YqNnuxSnVuK9/O27U
oWaAwsHsciBPbpG9N0xpo5lpzbb6EYKiRf+Gk+BmosQYtrBdS1g0IshvcuQ1fq965mX5mTzd3Sc5
AKKbj36za+WlXx04cmBQ892gt2oRN48cY8OLQU7BefxJJom+pWcw1mcYD20c/9zLjdtKYs/0EI/D
WiRDi3J92aaMmRoSDLkFhBSX9gWnRJDKe9VP6SvRzOMpaRz/YBAyoglWUo9xyg1RNbRKfg8kWKGY
ua3b1ltWgpsWONm120K+L2Ucpfk8uLiOYI2oTCa3KC218c2mH0dnQqAoExRZxXG5ClAZgTh9oL0z
bf+PzACVh/vi/S7/6xIFvO2u+9rrSXeIpzq2jzjxa9hEs9bGEkGcw3nokVYmB4EZGY4oZzQlOz3M
Q8ZbcvuCDG6K3bWvxlgZvXKVWC9saY6ZtOVpKG/WL2URl8+Dytod6ULq1+FG+8TY6OVtCjYYci99
1YHlC1QIQJzM4CbDHlGD50dawr3/a9neyjriqqk1OLbkNHCLm7kT0j0n9Ptja8isBvvg6sshc5ll
WfvDsqkI0K4wIa1dL0/eRofVtylRENJhfIUojZFPIexT67AJUBe3FgPzcfsOcpxcCFK8Bm2WJCW+
WrUeTbySFiUYAnZm0BSZ9CVy5AksKdqFwayduhpfqV7AAAImQe6XRJKislwk0zvp7jYjmiJNoH42
1/mCjKj3qHtmYxX3F4EZIWEJrHEU/FJRI02krRaTzrkeOO5HLNxmMq7CDiNYeeAheEtG1J/O1Pgy
4i2Rs+cwnxBLVD6N+I0CMtBqxz5ETwhn13fg+bswLfhBgQyKBrORNvmp8iyVXCumdr796A7bPCGK
KQ+x8RBIzyQ5ucAU2K+R8OWqW4v6BsqZc7LqsspHHQ0reIwt/9UT45qu9+V1tXleKULUijVIcTRa
y4QCkC0eNvyclG3CO2+hkSo4azvxc60rbQNlDrE21OtZGItPBA3Wt3lqiF8gFvoxSBU4t2KLtMh/
dHrw3cF622L8sin4UAUU5+JoTxWkkkkXfqPIXhyLvm31jZRWD5KEeqaMyQz8+DHNbE8ZDi83cAdX
0+KEW8rvbj9JWe+18OjRyoE0zXkiN1xEUFDdXXWnpLLC/G4lgooA8in9NTYBr2RC7YJ0RbxenoUo
sv05usTNz5aYypErjo6X2AM3R74nEVajI0mUsYuXxiNgb7CmZv3Bfb1dvQVJHQ6B04aqMiEMgV7X
9eNyjD9hAedFofo6Q81ZTVFKnIk+bNOwySRUMu1UKcz4DSCAXyguHCRwexrnVO6tp866geTJoPkz
6nhnvJGc6Gh/tKOo6iAcEWHDe+0E7BMAFOyq0iABj+jRdSxqAkNpgyicI1yeZKEHrGlRTAnbORqZ
Bu6n+9kaH2wLxXKl0XXuCOt1Hf+C7jwY5li5s3DqzzNDCI29ub2j5WC0s/qLPD5hSJ7OlKYYozTl
UxUBr4R2uzgFTm9w5FpNRWwgffncnXV3hN/gTt8bEqBab1G5lwOfhGSriAPY1k3wwr+wBVkmrzxV
KXjD8BMNzOJWXhD1jtyRIMPXhnG/o+isS59xKMaScFloPvrxEfh1w3tReAdkQOx3GstGJz+Rzew8
Hcw8lufh3NGb+26SPer6Ih6uetZJtvTORjA10zD3tcbCvgWDFZiSU/lwSyoTywBqeXXMPIVKXqwJ
BlgbjZhRwaH5VZcXotRzMOcRNJ7YI/OPhIWOnoXUEgLFGc34Ff4zc2A7Jqb3Yzqz1daDpLWYfDvO
Nxfckke+lwK/G2gavrQl/HAeVPFyiyWUK6okYrhhP+XMuHc73PwTUnjVaGPsPU7BH3LsZ5B5u8VQ
zcmdNCGhB5hh5HKqKWhAqEgRdL3M+38xMW1SIgeh9gQgwGvh8l2MdU+1b8pN27b6Ha81ZUAQyOqO
23c+cSEEWstzIEMkeqM6dnv5Iufzd2IQ5bTPK0XbqSMlpar6Q+D1BEuon/mIu8WPoLDcAQA4mssw
eBakEWmLQOM7sQej3smiu25Leyj7rKROylt9J89SFCk0GBtdND43ctTp0BSoF6b7h21hdJrlfDN/
dvsd/r7ts4QzMRH3+mo4ecZ9FrsqNXz0vBpqODsuikoOzo9KJnYdKRqYZftjZAE0XOj45jj5Ilgk
gd5/yw675BdvgmPCLL6S9+xzoAWu3sh31Z1I4HC/QR/tS415wTojnSERLvULlnob+Y3SrGbMhI/1
4D8x5i6m5v478TusRvsiWajCz7O7dn1GMWObSgNVPbKWuaOmwpwPJfCoTPcym+QLMOhA4PG2LEC/
lSWyJXWapa++4veoqZV4HEdjRu+PXCJcaWWoo162Sficn6t28rVoRwJGS6eBohLhiUASWvQ8Ikd0
nxbliOqtKBO7DHLlBBw71vowht2wEiwvEZDuYgqoZe721E0k6YcnfcyZ/crnnr+qsuTp7huDxZAN
tIDeq0FGJ7LCSplBPa6gupFSBLo3zsqGOh0K5fWfcs04/beuKXPKot8PeyOrSNvvIIyc4DqmgS5r
fuRp2NHX2bY6Sti/VErRE6Kqn80xJC3Jplls3XQV4JqU0xo20b2MKMMkXLB/SjNFFKo5/fTzgpGJ
jAuqwxjAN02SMAVxFh4XvSkAVt2LTcL8LEFV2nJb0P5JeVIq0rRm+3b+PZ3lUyhuK3V40q520yt3
nS6ZKOh5U8kgy0kxxRWZTzV/npVyDee3CmwH/JARkMX+Zl8gOk53DihRFyALLvb19B8p/S7ZuvZi
Szw56OJScbO7gu2B3Yyj2eUpSXTMRc094Nc7OC1pibLcog/kH2AuO0+sieBljYga3vO0zxwHnQ8Q
EMgPqtPtqkQo+hM8CIJCDRuh+zHdTym1AS/nHnVaqV0n7OIGifbIWbnsd2C0ww+zIlnnZjj9GK36
NRyl8SSb3n0wcAJjTtwao+ngKXiFvAlAp1vwEAL1GyxEpGoDb7ulqGbzdI6E1LCnICcEXmY1GckH
LjwaOsNHyMR3kCrGr5yIa5bNQecgmL05F3BY/I+Wz08Jx9GGpaTjAb0xKkwQBsy6Fshe0dX51wQe
7mbtT8eyW4eMc9x2FmNc7d6Gq+ajzHBzBjaoMpGyHub5GR3ujjQYrmWXESOn9yqVDEn6K2wGoudB
/zdkZv9MBvkpKGk9X5Ahnun5ZL/ZJ3Yd96sF7xQwyy9qlF6so3SHCljFyjgFQg7LVcCKdlntWVnX
jxFu6uoAk3a3ZIZJdo/1fnSOIqxTwPpr2blqzr0t0tVizG+9KFi3Kt6DcfJb0Osj7JISZVK6SDK5
16ss8bRjXq2BxeExmO7dOjZbATBBuh3WoVSYUAaFbMYVV5crcAhEvqNXg9Ni2ByqyHWf0Cg/OVJK
7Hy4mV9BFm/6h4NGRvbrjzM4/9qPiFPsQ9fHNf+IX4psZlmEY2eCA/bN/BblHWFLVX0amjpDzl6w
mkaO3pLJ9yixPMILkX5PQ32jKyYUJKSL/wDj6IOYOhFa7PdugM+IKLtr8L79xoAlX7KaZ5owHfb8
GW5L+M6G8P0yfnbUYaAF4D1teOPxq/ySw3R+mGP056G1o6fN5prq9bRTcH05pdLrJtLKWdsROXvV
kKDet5wkGpxqnsYBv1gNY7nXieU7EZfV7jRJXEzvI3aT7CY/fHMkwJmcEefc07tLe/hIlCdmONpe
yl1VlCN1QmgNKc4gJ9hrl2U5MlmKDxFqs9iED6PEKwMeoLe4h4tb8NOw+Z5F0OwyRqWgXuzXDikh
Fuc4PTzRPOGqLGEs8J0NDvn3sbaV2WOcszI9/LCWVr5koaypu2z9Bkpk93FPdpvOLkHsT4HGKOTv
P5AKfRYEGiOwnNGW9fEblMIpXmAs+y5pUr1fHSOgAmRU7M1Si0Jz1mobIstWHJm1rE6mqpmAEijT
P9Er2O/SmEo7ACccYPIEcW6aIiHVLazf7FBDgbEIYLV2tAvr+3A8/AI536g5oR1vq8tvHInwPWPM
j15RWAlS5ss15ChUGQWQQ3LHQSV3kJzuSZTj65woBOyAWFjJwaSO7r9EUvu6BDvg874Q0bhX2C1y
bE+v8FZAQNfulK82pqpj9C8fiUW9q+t3EV+A6PpJa3oIeMccfcikRKhIN9Byf3QH8k4bLlac9QIw
bA9TKr/ioz4SSic4oOaPVqU3C/Zww49Tdfo6bo58j9G91Zf2V1Y+3t42wMHjkEuLc2maUfoCidHz
OYjwLfLzuhysl4TvFSS5E7aO+XSsJ5/WglJcZXM5nGLJzjmSCV4dqLXbghsaouavGL1WtpvEnRSH
Di3XAMcn8LBb6n0J5lpR/rYMz78xM2fx3EutGRosxqurKYjLf/OMHVGktzgwG22znd019R/j/WEY
IRoMMe5uRbxGXERJor78z5kcRRd5hBBbPLSxaFYFBKCjxPzukKSPchk27nas58D1pPpoSFc2XEex
OvyCbmJeHEBsolD2JA3k2rWR0hdmD2PlwVYBNqAv9TKdHLlkbcn1L8d+Y8OF3McARfQYsn8D966T
aUw7WFQ3f4MX4efkr0rVQaNP9w0fQAqJmLSC2J/eE6PVxzr7Q6lx/0aEUGJdQPKEbvLH/3bFkulR
ZXhrTeoh1xJMJa8d21RrHA/h53Q8JGL0EIHYWtfI8C4QKzHMQKrZNF8IOdZBD63y/2aRaQzr5glb
IH9kAy+W97vExTs0tNn29VYPOT3cNhk9AkWNF58iDUku1Thl1/bdtisZljh6bXQBHlBMUl7DHG3g
HRJC5XOoJOJNd1jIbJqjcHvk+dpdgs44wiRyM7KU0Y72EkreQz9ZB1Mw2JhuEhJbvgCP0rsdZhzk
7a/srOkYRTVji9cGAtv/YhgTFE7TaZEBue4Zmh67rt0fqw5sZ9Tj7nsUawOMh03SRVxvc4IAg93M
41IDk2HmVi/r+t7713kP9dj1qv3XE0D/+fmxyqzk9tsgBn1VHWHGn8DkDLixZ2e7k4hJTdckKdfu
M1WuaMIXpCRpUQDiCSQTTTKcHR7lRWvOsDwbuNqHc+++Ap029jzYwiOFX1HZ/hqrNJmkeLdLKSiY
0bS4hUHMK5nULMc21lMyzOf17pneGHYPHkl+l2YYPuwcMXaYM1vaXGVqTHZpZc4dyGp+yi31mqEz
NiRsZaI3a9GCTYOYoe1YDKTBm9xSDlyqbH/Fk6qV64M0GyRTO4VBVD05F/f7U96uesWn8UlJAdFU
RgJxxrppU5e0eEiLSYqCes5qRqyOTA6/dIJ+RmZ+Xuoxb5aDVlpv+cP0TEDnGgSFyQHFwHXOkOrc
HKwgz7/h4vdZv2Orrj8uynSq2lVxDllZoBIpypNngKcDXvVK3Sh/8OWv8rOgEcFI7BJs/J86ZDeS
5bPthmVP2HhkzIEp0myY+0Za591HZEAQQcy5+AdXMl24kQrVp4kNFsD4x8FcAd2iG9/5fJKKvR0h
YR3vJoO9BBzuDxya6tXANAFSSnotMqd+kWKnqi3cx6fLlJTM7cqKzS4NJJbAPjOdtav/7GGy4KdW
O/JY3W2/H24JJvUbolghmFvEr+E6PdTT74GCK3vrCMIzN7vpBjTlUVOJp/8jO9teA7juhOy9fK9m
slkCRWJZIxVN9csBg8RcKYFCYXXhUAO+LHcUxdMvYQQepzaRGtGabQW9TnoBVwvGGPOGmvWFjtI+
Tvu5JecePyAJFJWxCa6UAYCsj9h5tmtdAvtpZ9uXBVfnY1JJgOf49IelP6eiGEQUuumTKqqf7VDv
TNHZmmAI1mdPmnCLYpdSCWr+jYgkvj65WKmkK/hw4MkzvdeOHSqJz9sUZZuNKSI+sVdGJ7st1CkS
ZN1H0aVtC3YG2bqXWUBG3rIuOQ5iz30bp7av7Oa1mjCcfQ5d8r+cR74tuv1zjDB9Q3XaIUjBpm5S
BE1cjfVTUj40oQehIR1bcEIIMjvzUpYEW46YVzFnaUyEMT44azR0WPBbWQeo4cF3oNnDRYISs3Yg
8AJRAJwJE5HcSEiODqWJef77+oV8sYKZXlnq15tkJ/RolYO4ThJFTddWj/BJ6dEfX42z0gd5wcys
k5R9lezR5JF45HLGv4qJxxyY94jlUZfYWrwpamnLmiXOeoNBXR22tNtU0drYXsNtqzkzr3Kg2AqV
bxvT+3pGQXMDry+UeNxTHAjc/jEB70G6iERXUhg1AH227KuaYCGCU0lZbeQgtJduHeI/3lP8umSG
L+dVIR2WjEYiYdqNjt5De9BqyLM0AfpJ2vBGQhsx/f3nCQaFstu7idI5dmvzrvsBiuGybkhCDq1+
8eLPArJiIc8sjoanMBxITA61CPFUb9xFiWp3uUIG7fWZMY5nuwLF5OXoX8X7JpG1UWIVQfAqnjoF
1E7wicgT77BwI+4MK4Ucs9Xb3xDh/0hAvhfIZtFaAvoYKRYCfMbcESveeM2or8vMeA2lVjM21G3B
mhCbxHJ28X6mLG25Ka66qi/TZb5I5vxxWj23uzzCaREnpwRQl1u7kpZyRQgvUWdzs7SvxCpJG4FE
WBjkRd8BO7Rb7ganqP9am3ChwI0b0MMA4GfCK4N6AqUi8tAsMpJLnYPUpdOCdlNKOtAEE5XTGfag
hl8/E2pmoZ88wK+wSn9vuK/Kiak9URXoTU7ekeRj3s8BKSU9KrOZTYTsLvfUyNTaNqFM4SaEtVgK
c6Yv+wZPUhh9LKVs8to0ZX806XZUwvq+An/8mjboXS5t1SA21Mh95kQQO6WS2Lv3Aae7pSrIWG/q
xj8u6EyFQcsnwBbzncF3tD7oB53ErZsRvA9Y1+DkXN6ztY5FjTpQbbMU879aMB2CGvqhDUTeebrr
bwTO/4efGhS9KcyhNhnAk2Bw75WuCFE6LpOPJ86+PzrsDjWSEDF3bgwg9x08P0FX6O64WkqHvw4f
QfDYBtNKfiJOSj9Kl9EXMkkAVVxiv25IjNQOhF9drUvDjg80+OMfHGg/d60gpZrJy9t+lmlSid46
nO8po5fub19boklDvA/4EgPBbGX4YVFp2wy7Q9kyREaUECYh+88zZ1S0tn8fsrZrAnDQd5N6kvP8
0hPtfukmLSvDFtOoshwBYV9denNxPq8Dy/NdG+r0xVdZL+/UqTxhG3H8ac1sFDJGEq0g2RsNl/5a
P/1kg7wUKPslEEqPqZQaYYrweCWxv4RgBP699Twri8+OW4MSCJxhxEhC/khHRYQLcgaXuVXjd2yz
lObWSHtn1i9GuwBKFYeYX0urKAuR9JV7II8C/e5tVRiJ1ikHsu0b4syqhV7RvinvxK2xMVPYFPyd
iGkxvmzMlB5TYA32u87ZJSvxi8pgpe52Rof+yN0eQOcUqrb2ziUq+ma408wemkLHMS/hGHegpQh2
dcthlWZ8xC57J4pbR74a6cxUp71qEvMb6MrvME8/NBxvdDPpNZy6iawryx0PyoNJPnRDo7ZEcycD
XFF7NzpJD5i2yjKcbs6tuACibRKDmkytkQeuRsnaqSVVAeiSpwLvJT4uYEKPNTJ3sYfLBohzDc3g
pSVUcfw+VcKdn3U5Vng0UzJ/EtTTDQzWVyCu3W79qYcO/XG0hHn6jO4JEpb7bjU5UirBIW6PLWP4
I/VZFkJ6e8l+eC4tYYoM1HQUTx7vc9Ku+7JM2bvoeIitGCrTo/I0AIlITzRnIlWK8uJJOrelEqy8
lTDNTMtC6Gx3RXU1wrvycN1j2AnhPNwWCnOsm+cZ9DLVIabt2JtJRp093hI+EfqUME0fCxzOZOKA
ncg8iRDfUiDeLrTlUE8v3Ui+XrAdBrR5wrHzt+XhmrPA85nF1bs9hj6MjtC835683YqQzD3/VPEq
hUE3EtRyzF7YNhdZ+xXSDG6j32yMAp2OnmRD2+50YgCDo+FYXwymAutymfZsxStqcAgbGjkgRotG
Axlurt+GBfLOd6mNo7ot6emEI1rQ6aXaDrPO914FUbtYczUoAvWA+wpko13BFlHKORt4uVipgYdR
gZeTLf9EjD0sqHae8yVJvTnCkA+Q0Ov2crcSzxs7hWZPY3wdjTZCLIBs0l559yMtPFjmRLXio5Pu
xtC3PGnX6p5i++Ik9l3XxxZ2MtH7U9rrzQba11wQA4KyqRUgvekzW3rw85ItrruVob7joyeN4QeD
QMDuonW15IHeDXkv4g6JGS9hzQTOXRzJwfGUIqD4gVz+/AMcM9gbMy2aRQ27/TwmR87IRSGyFLB/
0q9QZf0KEOCMQQwxQFfaiPUUwgRScU2Cpuv9LkgZy9VCX79Ib8f9aEWXYqgKu5MCF2UJp8tdXXUn
lnj59uZ/Vch/5KpB8isg0pigyYmw0XOssi/eo6xMnZmTHDeEorQnz/PkUkbqOmJhNmKGpXZthqGu
t89ZFE2lvvtprAt93qBJja4pULRg6ic7odXEX6PeBalrFaiQ3QYWqwzI5COCZy7AQWiQJ/MFa/XU
F7HxL0gZM3KyHCSTTBJ0T/FYNqx4bRQjDjg3qCFtkCbb5+TBRFEufJ2jw663qC+LuS8yGNjmRLHg
3JwGbBHg53sElvGssYYj9sqFo3Ee//qA1OX1unc/W/UFDeUuM+ds/9mokeZNJcoJumS1Im7qm8ns
b9wKjFnUJMCyGD4Hu12ZzS4LtrFRbK6Y9VzybEc/nW4Uct+29FQAGN8y+NFaJc7vvQBa7jyvOiqh
IpApwjcwdXhY1MYshmedkdH4Xt8MdQbOPiJ9n8gr2OMgArksnSvLLJAm6/zlIrF7UI2BPywEi2bZ
89LzH7+sNSifwbxeML223ebgJwBcc9GCSW03W5/pzupsVVG3D1gG2l3H9OEWZiEqW+D+AQDTy/mL
q65xGki+gk4t8vDI1IK4uItBFyKw5pE4M4ffJmk/RGGYrAwKQFXDqRVrdRkDcVzq58DRb7H59sta
HknDgsdpM8BRz3fUVgnMUG5XcHWGNdMuc+7rhEv9zOdiqnDaMS3YbqVgfTQOr6RQMjaiWtTccd0W
TcmZQ7/9/zFns9T+U7jEWNzDVNn/vNiLcpRM9v28xIeB2xAxGxl3P9FgdzUySYKrBxZzZkuiH1Ge
wtsg95MOxCjFofLT4tHZQH1zuACmuY4Quv/wFHorbXUMHHugnMoFycHzWO4FUCSNi869OniA3nXA
/DsKWDjGphN/Kppu5laW8oRQm9jbR54MvrJgazADQTZo9XTy9Je6OrbbzvUyKgFpUV8YUUpLOJub
vdnAl5xDyBqkYjSJiARLehL7vyV7A5VoGFeaJ4Tsla9XZe6B6B1vSHD/4nFNI5PsuC80AAJSWeyB
KaVhJR9A/Oh/s7NQrihgIZj3mK/3Cuy+2OPPU3awmv+jt6NGc9xrqZjf1oQU5aZLhjEOAA6tco/H
PPg1L/BGrCfVV3JbpQfozczsRl9ga0L8w8znVLSc9/Fvy8YFfTS5PKm7iYfZwzjVIohXKS4ULSe+
VKIrx+aGcWVvnxH4/G+m8ZNY8I3jxF6+N3RllqeGqPLn9cgo+wd4e3I4YnH8YYgP/eOZdjMXClru
d7Wa8023aSndTjmtf8kCEfzcINiIycb9Rz9Xs3LVhUoHpuDzZCRYwUac+2TwVZr+utL5da2aSt1t
C8V/JVCcb0MRoK/2zZQWDhjdw6fvPXloXcuYLL8+GmRILYHoXy1aoPbBXp5D6yp46li8W1WmyESg
31L14ywWg4InTRNZ+m7eNUZVm6COPQm2ry/FLJgcYM3qSp6dYkvCGWjIGAkYAm1VcyWWcH+EIojr
3v/742XtF1UWnFh5oWHqhe7g+igee1f0BOn4Zfli+U7kqFuLu8nzdcWDWJd5YfjFdzfchT8V7jya
0zRQblzZi8S3FKl0sx7zodUGL4V4/F5dbbyzyRVN0ggo2nDBGGP07At7aZS39apjL3Vavku1Lg1W
BhNYG2QZwEM9Q3UoB2WbwyAZh1FY9KxEcs5lCyupNJTnOrIAUGTbtGaLvEEYh0U28pHJwCZD6Nq2
goV+f+UAMJhmjtgW89G0GroXZxPoNCbxNI+MtNYXA1M/lLqIKkK0DkBx2ztiGjU2j9l0FRJ4/gbe
3STeTKbk3ApoPGN8p6cgbTWaxwh8uVaCfTA6vwIxe25nyhAwJ+TZCBABCpYO2PyPgxqTuEKs6EfJ
H8jLPnxaCgwsyQOrawCdsEmbBG8nzJvJuuFA/3/837lIs5C59BKkDsui0ytaTEIk6ceQ1QI38Tso
JQYWQp8EELGLw7QsOP1ZkB40VEN+LSGODFg0VG9/MyQo7cIJH+41M45EdmOU74gOQ9QSw3SPXO6n
00XtKT37YE7RTNmkTpzUSm123WgCL1vK37/dHSEPGow0XChImDEcSPUL3IbGBa/x5GQKFMpjQr+H
QoYUq0CBdiMTYDnScxVduNzHNaokJ3QbX2njFIxSfPgYOAoHbFGVpDPvuU5hOJmRyZM81UAZVKzZ
ejNr6dXqk+imiYTt3vhNh44UWotCelcQ+0yGarORGHEgcVRz6mTc5pVc7eQkGcsz+6hZKFTcyDpv
CLX5OQntOqLk4AhvZ8hRVEnVclJecztVbB/5EAh/4pRvxHJzwXwOLzTH975uCUOzdTHaGVaDKvf0
vYzDTAwJVmp3NbdfgG7CYsaKiFVNFKBJkA55QDlA8zs36JbfZ0VHT0VAxjwm7RSrhTGLGFfIX7v1
zX8EEgBMxWkrl6k3IRwscboWleDMTsatZVWjihiiNibaY4Djyo1WAod+FtX+B5qr+B5XtYvZOk/x
kFV2e/m5Lq2VW9fJKA82/XasybDaZoXLZOX1CoweizXXXWGzw4Eh1uDPgw5n1VP+zxjjn6y8Rmox
BkYMCElq7Rpq3s/1UEpCdoivXURRS4tBQaI22BnOjRQPG/C0DVrhhkK7l0jy6j+5gw+RVz8Rcq1w
/ePVXsT6FzdB90S4wg7kQpKeS69Ls3VQqH4Ln7B6SidXWZgN5fg/3aMr0rKOz8f517YO7opY33Js
NTMi+f/6SFnk9eil6AOUD1/2+p2l9LqYyxgTI3HGmpSn+/VpumHBRw9NF7+TnqwzAqoOzJ8ddIVQ
gTFy4+4bcVRsjN5WU9wKT1xgOsLHKs+NM9WAbneFwo3FFNXMIZgTTl69qaA/hFkAW8hAxAIOfkPg
+nQrWmvuJGWINDo2avfvjU5420IR/stcFsr7IdQKe31IVcxcHjaS/dwVHASREWbipNvLXMH+NIE7
5BNJphgtYmEPAl6JbeKlqBiCfQRKK5ocy4isqnACamagFJNvl4IDrUr2mX+NMnEjm04wZHQrdcmt
re1BvbFldAKQQ5iApAlrkD9exMScJLGIt35mnyyyoXKdUqeVl4Y0aIzNPBoqQX6wm8aaazfm1LgP
dxfaPtANMIW4kDoT0SPBRRF4naWOU5QCkYPtBYbQhoGj1SPy79rH82OP0sPK7PEUXm4OjxtoSbTl
e5nlbWHq/ZNc1fPHxJ2xufft8XwN759e7tVPlXj0iD8FiHbjYyHnIWtSGww0RMPyA7ZV997aO88Q
wWh/p8Bci66tn3T3qz0h5CpJpjckhAZ/kzl4GzW2TH5VoTv8+XXWoYEXs5obawtcXMeIn6XsGQrm
k2nuAfIskSV9Nb701+kO0giGWzL4EdvVfXZPzgjX0QqVe/QbtwXqw1dPCTNRlF2o/Ym+WZAHd1Ox
AwyjNbl2p3XpDNz4n0boE0di6JpSmjmpPdo+qQBZny/sknmn8qMu/ktVqizoSpjPOPN/QmJsaYDL
EyP7c0UhRgrVGl5ZBdUnu7BxA5I2cU2W1LKGKamz7ByucAQeWUIL4Kol1HyjIAldtVWN2K/cUZYe
VH0gSWtkRvqsFZdvWa/DOMqHhguYSg6YkwAvOm6GldpaXyrVj0as9WTFQaQ4vlzvBnZBiESFDjIm
KDEbt4CO4AB6ywNtqKZC068JPixO1yZQRIBh9MTrvIsDMt6xRyf0TH8IwlSbZk2n6YCQmYzsVKBW
YyVQa8XWv10FBu5m9zxemf7906LoPSkfe2utN8SZ6GZksf5huhvuBHia20Mg0dHvU7wQbj9I+Yf/
wWoTSdXKYRL8rA+DJmds0r1sBYDOQZbWoeObYkaymA5AEUK8XiBXYwMQwFdyTUA0U82mC6ybjkjz
rIlhlJHldLD42qpyhT0PYtgU8uUhJx5OvLdpS0+k/EZQvaPBgkuhJh5ql5SI/BqjWHdc5ik3HHPD
6/ggilhrIzIQcLBAbDlatyALjsa205yc4xrqcWbNtTAva2I7fLIjrruMoogGAOtLyN4nSfbkBHMp
kTJZVRERSKrjVxD6d1gFAGluDOCD7vbZkmT6uH6NJZqU3M/JM0QrXvTA9TNgWfdaqUPCv3fLKwiT
o52y3HyyEkJvHmFIIQra0JRi+eRqse8Kd8Dju4ve67Hh/hSa9DmoTYdBHTwfknZGY+L77rdwwpkV
/UCEJdJimWMRZl+cwz2+fvtR3Ywxy+63Yf/H91b2djC0bGA53CZxZjknHUYc9BT8KLE55JN1e6zY
CiCzuRVQoNkofsDomx5x1rG6OY8nCjvXnIkURuyBq6Jvo4Zn4+InZ82YNZydG5GVbkFwqqSg1a+4
6mq5u6ErpZGJ+z1sDnzzvw2svlcaNAFQukorlaV5ESSsjfPbWttdkCEkHqmQ8qdJaecWV6jnQUQ1
ZIEN9nCOUIuJ9IEgppleV2Plm9OQ6qPhm6RDfQshVGT48uo2XBJ15nIDUDy+z4BjGysuMrIZBBmy
514airhjIn1uiiq5qtOSc/mqSuDwAmQIa/m2fCLjdYNClz8BJUZwBzpBKOx4drwX0z39iClXo5jm
SJpJba1P5w0Ng8VGxfZ/et7uVZbAZ3BV5HWXt9m1uEqMImhvcGJMt9cUf7idgnGS3dGfb/XVUly0
vWcH97eO9miCKA2m4EbFd5f+aIcrSxBHuatRXudol/3rs1Y4QUZS0eCYkkJhC3dVI3eFIK9PNHDV
3VGYAyD+sAJmdU11ZtUt7vL/sIEpANJgyA2eEMTY75swS6GUcPQMVsMhQJA6DGQNkbaB86/8r0VX
LoKb1orvpJmZ0+1aHxLKHIDWqAmHosyU6NTgwFOlKCAdPwWFiXEsJIyDeYI3BS6FxSvHWotd5as6
f9nShXWqBDKpxro/r6MvVtQnUt8sT744rrqNkUYHzITRCSCXgPOdRnf8felRdGA/YssKtCLXY2nI
GPZZHawJKPJ3wHdQDbfrwJKubl0nt+WxaQ3vXrLFKXi/bhIoWMxG49t8SbOdcfMwMm3RatED4KVB
4WK/FQhN9b95D1P36qXf3FcqZdC23AH0WXID1etJXpSVNFLRW2rowM5xG/zQMflVm9GUbk1fntVz
4su8h6F6iU6rj2Xfv4kO/lCjSWSTnLQ827h7AEz1pQg4Pb8i/zc6aDWM1MV3dd7Wod8dLtp+MOgm
SYH82UnNkTIqIYCWouuZiDmJ1q8guXZdJPqv6p1+mKPji+HEnyBHsv3f0NHO3efQlScBNxly5De2
OUBoYLKUQDjwZghRK4p1gTR5QGwtfP72Vz8YKqhOjWBZhgDLUTZw35GdHacc/mef1Pk4bonnRhy7
RAUCe5lVxo16fnpL8f2COmdrrTOBYJPRbHqobRVYJaCI5tFcbFNHWoLlEj5Zo+7LTA9GIuOdqwAB
JMRn62vHlVjO5JeyQ3M6N9YOzRPXt7dlKIXKG8zRlNdMtzKOBKFmgPZCWblXbvavE21H3841IfZh
7839zHGBAaQaUwxiNYV3QJo49WbnnTED1E4I0qmLXCgAMW1/1+w96FQg0ewkrBpm05SqrAOcJ3WZ
lZ4vLtaTvwlms1o/Oq6GjDiuEiEmOS2duB7o5iJ80mk9Rp14f1v56qfdnqdQL/RYZb4rCmDsGgnF
o8bzIArQ+Qe3aUGhCdMI6uu9ZXrmm27z1CDUHqKMw7kPcyUxktAX9yn45g+ULbiMYlz82BLuQ0Vh
bt0TRgnohprW0wXK2IKZ2qPMRDxOlelgDKj3bk/5vXQzgeInP0+/TrHBlumruduueBbPitisrxro
Pp25GI01O/gHOzKkyNBa2N7Oa3g4ucvrMCSxfAmTY5xy7gupgTCPFjNtC4t3AOUNFrX/I24Knuwz
NLDgKQzDCpxAnqZjhqNEynimRRpFkf2hReMmvg7k1edBwKui5X4PHFh0ICdu6q1GbI+NiKFPcXXq
sd6UXFF7dthesAvmNBtc7jm7p0mOjaKuNEvSx0gTvkS6U3+xhFdtHLJmzgMgphdKe+fDXjgVFtQo
eO2RH8G0ctPIt8t59QT3Ie+p/j7egp6ZONYJGgj5HfI+iC6R5XymFWKMW6JrzaT8uQQMsKe9/Rba
IVyuI48WcYj4ZCHZwjxxLYEfGzXJzA7E1cF3vF4MZuJd+4YjJbj8EXJmAj9Ir8CrTICuqMDGjaME
KXPraw24PTdseQdVPFlqEZXRcZPn2GJBTAlMqFpDRhROwUPNmWAFfLROZiEnRHulfzLu9b/PonPG
jFIB3T3LdlpOA1qwq3SmUwV0TFIpQY/IWK8dAq3IfWCO2Owacs/fOkID34YcOSohfnZaxPYRb+JX
KPZuXsI1DdhT+wC7gBZ0rVSp98GLIPVdVVJv3IcrOTu/E1rOWh/ie20xbc8Wq2M1Pac1FsP/CFiD
JAPkMNB5uYrE8ONSC/YPZr30g0oRv8xOU5Jsx5fuENtcGmJgmsFERRaDkQegKXkiq7M2QJ+8f74W
ignfWCqUdPHJdtFVYdR1X6Nw2p21hCe4pP9LW72QeqXMt8t+IsPHMZVGzoayi2fJw7ci1wBEonwD
Q/9pbB7Y7RhkwoKol2Q1j8Prj5NxDkerumDOBSgGHsGg+bpmeLZDg7mO3J6SfzdUMNAdDhDlPsiJ
Shd5DXTh08tu32Fv6mL2Q0hRjEUz6t0eOUox1sWX8MeyC7E/+mNgOqyHW9uEedDXUgEPAFuWtjUA
qawdESrqldSwF2zHbsUzyGPWcEK+Yf2QraZ2+oB/BZjp6JtigoZULCDLdDsxeDHH52puCnCPWjoB
S/1nWA36e34YpkcIXGj9IuOYGlJV1izh9DxjuUy4DhwZZB/eVxNFvjzMsDjTasgbqSHJhOPZ5Gds
eqAwngyBmHkpUw01YiBqp4ksrP/I6/8QXATaeVZnUMG0pU/KQdS6zS7X68nziSRrAFvmVkdJ5mqR
DOaU+/BPM+Gf9ink/7u7NzmWswmoFcFYga+O8jCl2iLT/jAgzODWEQ+Kl2ZaIQe1xvyqahV/M2LI
oYKAVL8ZoXQrBO3iXjhQBNRQlzZarBf4E1Xs0GfRWFkeJxShFyFEc9b8r9TVqGC0xn63/3gcR1yo
6aUeI5tW8YzbwbfNOGqoVO9rf6peXX0BAuustkJ9WVhY/ssGDj1jXQWa22x/Sigr3jkOvqXCfLHD
hT2RbjJYeYrd4xTIhHOS0aGq9bt3q/l7zrezZtM7i//XllaOv6mY2TkcF9EpZszzdnsEQedns/YN
EuhjyvL8++aEsj8AV9ZIY3UVTMlpbpBzHfXZNH0VLF2xe09aKKFMkHyeJT7a64/UTfJHIiLlGZPG
1l9In3YjpN8RH9r0Flts9MQ5ArAVH7ExpW501b5NVAB4R6Z3U8JzfI5gipFG4Iztadg8mxbhHlA+
ialXviKCT1BSKVhpwQJLAWsM66TelHy3CvGiAqY8Sf8Ir21p7qmsck0Sq8Hwgab7PPEMLmI8edNR
kpliye/wS8Pc5yCtcqYCRGobwGWWSqnEF9OpPwuWVaTPxflUmIgxkxB1AUnvWupoWqadXfaYuF/R
rusT7LFhssR7iUhIGUmnHwgy7mkXccwU/TYmAtgzTTkeK/1JZeiTlL8ieaXvrJ4Wd99hD5bICB1W
dRlQjzPr/LF8NQ6ZhKKQ5N/wiFyEpgpkX7oC681M0am48kQ1xkelY+eL+A/qXY/XkoHGEKRPuH3V
PMgNZtQy7NlF3/9qCFi2rKQg8x/dIaXA0DfCVvMYhG5c5OgHlnOjzwRydkZ9tLOc8lzMcR4GVi7b
ggaO+Ac7ok6//Sz0+uInmvgD6TvOvliOJ+ASZb0dPZvoeUFI0F2+/HOZjCr0RamZ5UhUn3egVhL1
cUurhzNF1+fNegR9CcFSmq6TwPf0gqZH8qye2Wg43YnSwsWzbl4FKMRLGwFAujDLOoyWzp5x6QUE
8mPBsNAhAfsVJlpda/yu9CaUin9mfuR9yVXtOcnEBWWvTSnPimWE4VHAYSjk4+9f5nPd8JYuQsoH
vIwgEaga6Ynjyh2U67ify1YyuV1X699PDiWDLzMPR0a+buJHFumA0TtZfEaxUC960/yH4GzxpVUk
nZwGd61L+l4N/iMolwaLYowTCb2ibDgAO+6iL3cYYbN633wmoxYIaPK9aLOu25NH+mkhQUkWF/Le
jsX9SQ270sPM3ee8NQvJvkNnGVy9nrNdXBpsQAn+vwUiNllALO0xFgdSLxkQv+ST3/nNzUNI+UjH
sH1jUnsGaU8WzugAqrm/KvAU1QlzXWpCm32zWfuCrakjbECBQMMfhAJ+qHN/HNHrqbBYFrOHvGZo
p4pdGQcCwVpFSVFRPMld/T7ZpwR8fYSz1LfcXEKkzj0Z0Kh1ZRjehsQOYMUPRR0Qw1X4g9P6gcmt
AoFv2vH7s4CZg9OI03ae7g4nYVUFxuPCJTOpNxR/zbkbkM25o6/VzJyoJpf4Qeizo2gOzJUixMih
CdlT4Hz7ItuGP6/esXp65rwAguwIKRJQkS4hP9u9bc3WtWB0hnLYeNYyG2Lya8/wfETZpvkA+DsT
FIXMcP8AIx6fFOUtsizZnQgYHhN+KE3/sMvvqGQa6sZBpS/LQu++JdHDQ0Ma+ZdR7sRPNTtMdFCV
WUpXfM2qMVOpgcu7fuq6t4gPziPw+ToqyAz6wVimTTJdoX7EKXBMsI45hGVza8/FWmB82ROteThT
edBtBkC96QcRQ605NidoPavJuA8xiCqdQbL3Eszo+2H4sLzHZGKQAoxs0cv5ChmLRiPaxfET/NsI
4QhKCkt8bjnvj4TzweljsG3jP9lx5x4zZj0RRBeGqmCwMYzMMJtMnEEbzb/V6FqeihuX6lyqjXSd
UslHKm6QjvTh6LdpPPrcGWYStKOSc3oDZXhoVzoEUIXrHq/V/lBcQMvteVs1hzvq259yMNIB6uLG
LxAcNLX/OyKVXlx7HGDHXXe84v0QjJrwE5K1oUaMxtfmRchiy4VtjVDZFhErtHgF7rgW0QkQ3Jcm
26OCbpndvO3OFseWQH82NHHCdrxE0nUtpFbEP4SC4VqW6HiD+LjKucS3zX57tURk1heE6xw5TtpX
jGJr1c9xzlaEKw4aBfgo548/4ofXxcMs3wtluS6RWbJUDv1RLpfJege1D7i6UOp6ueGopeODLMjt
ZDFzQyp/XxvDbw7IxsXyeXQO907qntgWV/DL59MWZ8z2kSWx4HcgyS13oCE3iASOb8aHVQ3Lt7bc
95xACMVgamGOoFDU5xkWm7D4iRsfToxlnaUlg5Qbg0PUItaOgqPoH2KLkjAhRGg9O1jUuXbCSJfo
7t+/b8Sa/JaGO2a9+6wY7E+pu02F3gtejfdZ3esl4k35L1XL5OWgCwlwfUStdJnEU687n2MJUp9O
iJ3ufRoJXEBkkdI+5daPtFnLVnw8zod06wilIjWrtxw1cgBhrR6Hjg6ncfUZ+B9hnkpGqvai7QCc
4Jf+2J/KLUVDog+1aQJ2mU8MDtmXO2cJfa0U3EOqgdyqa7cJVkL1huEXOmBLNb9rzkjqJfmWsrJl
xIrhNEXvi0X5sZX5MOChn41tWRPJ6BOqMqL5c7vxNP9adkSeihCEot8RJQ1JIOmAO6kFPG2eAr5N
qDMWyMBPJgUkGFeIS+JlAeLhi/USMkq6/XT0H04lVWSCU9t3+nha3DFwt+6bX1RTZbp1nImpQZs7
w8+sH47hqRr7GqokeH7vFy067K4aziNKD7DPLm00OEy7P5irrVweLSOXyLNXM1p8ucGcxvFMVbk/
TG/tSUhUVDTXhWayJbm00HotIXJRP+45O5WJetLVX7sMPWT+ZGnkO3+aDuSB/NHu4VwOKT6g2HiO
svHfQ29M+LpYWldE7JhI4oF6JzkP/SM+PPvdvHpej2paLKoKkpZZ07cddvsylU5uDIFWgztcjtqQ
k01IS5hJREC5yTpZjV8TV3Y4Lw+vLZjrboEN46QyfooRXxE8bnJDAfhKnsNKOsyPiJmYRSFAer9Z
N7UYPtDw3RFtzvS0M1PKPz8VCifHkb9CswSPsmW7JrU8i8Na+B7Anu6KhRTKmaQh8stfxyb1t9RC
dkVWcrLRiXGFYtuzbCwuK7XLa+yuaYorg2M1hg8p6BMUJqxwOaoj3dhoUDK3ubcgixCGzEau6wng
evgBZohduvZEIDO0EKA6EEZxJdNKAxZAPOvi4bn9//Kc2l442PsTDVNTP1iZHwnjWZjioIWHlKFd
hWTjc7f2VAUY0sHVww4NwCP1fD38/wOjss/TuH+XgILDOAMgTiFl6FWxGT/HTWxAUfxpNKEDQkGI
fXzGl554GZB6/5311MGrW9kZm9EBvZJ9/gVEcAij6GxvIHMroUf/VCnzHx8McYa7gqnZo7yEu40T
O1msngQoZHcn3g/HaDP3gtIt5J+mxjKvn2Oz5uwrrq4T7eo6hlVGep997h0Zdi5mQFsz/iG1rro1
eco+7+4tYrzgRpo6X8weU+AB5O5s0gqSW6yCS1lbzGZnibZ/RBuupJ7gyYcES8LQVlUDZU5pHzhf
zsuNjKREWSG6ch1TtJ/NhdfwvGVRmyqE2WqcglFj6SQDa3RqPeKD81pQoI4R31YE4hlT7Y1hUniO
uLD5j9MNIdwz/XvS1Oce7m2sDPVtrZsVY/Tm7qK0KGsRnnV+vPo1hB9e+wrjxnVzuZl26dEwtSJh
HBFCoTU2YlXLsS4PsfdRj2ndDJ6BcxXUEQEQ79GRorZtv2eS5jUYHDiBpOZxZMAHgN0D0m4u7Z3L
CSd6vsmdLROsGRp/VLZ2jmj6OAgPCVvqLB/YHCMlc3ztOiommBEOlUCvprI7MhvT0riLqyI2AIk8
xH/eX+vdydrrmjIDB5/ZPBSWgOBQlXkT/hNc9DE3Eqcw2HYJ8LsUsLObTwD+bej6grCiPbuEqbZ2
FNxsBbHjiVJdtTH7b6bgZk2HxURzVk5beXmhV8Fcpx7Z3r1cGC0ITUY/9PbicMNBQNInMIHOXFOO
vab3Kpf+oNAU6hLl1TBOxIXgRjwoN4lTSM176TZEIgeD6JC5XoeCwYS5Jj/zE2vOXiwPvhHqlqgm
eG6jyxxF4tZi7ZzFZH2ONOIpoKtcDHIfVO1lVREd8R+LNJMpm6ARADdiUeP8xuet7vK5WZbBrkLn
qcnmzXkWqEP0BItHb9DOCi1K3BxTKkmErDVtwQwn9b07HV+B7BkMFS6OfpTZpyfzlTDj9a8ozPiK
xPGzr/ulu3KNEBYplhrSWqEalGyg1KgM/xGw+Ts+KZDvnftbfHKibK85FIIdgxcoGsuE6M6x4A+k
8FPYiOJ3cqtLHATpyoJ04mLj5NeBtWwf1Y1Mgh6fyCF7RpEwxjhB2hn1AN6r+V9iFTH0T3X5DtiB
yEMbfbrpPR4PsR1wmn6V2jSaJ8wUFd6YnlujyYmpvtD9rMpTb2FwLdLy0NmEmqgqKbc4f4+V97K5
9MXk29jH73YC8nAkHg+aw+SM0ngMy6Zdm9LFEDgIUTlEefpGgqZb9Wy6LcZsxF1FltT/QU1adkH7
AMXuFBvf6R8qaIKl5PAjA/lSRRIUIzhKCoDtYlFsE/vVrilPlqFOZiowa7A5e9uy4TMD8l+r3IJD
EYw2ID3WZubBLcI82M33KmMF+kercziod3c8bAWTtC4K35W6si6QSjEqYu2wK8ZB8DmB2LVrvTiA
uLWPmWDzmAqWfjgaMUAwL7b7o01FEj4AjJD3bqTbsDUI5L8YhgNgvDZGTTaO3h8VSjZFQ60+FoJe
2WjFKKPF0a8hmbPthhcxmMXZLSSq50h+8G90lerbn+uDwzvt9NsK/nb3Hvrh4nKelsiZEWoajiNk
kIVE7lXAUvAJr1wZIjVYnrRPa4GuNrpfGKznwogN8ETBEttXXR/dlOXnaZff2/TIVB7pyAmPmig0
u0o5KrpqngtxBnkpgLzcshNTqb1huNHrw1T0htav2dvGEaq+H4euamFzAcyW6Eb4/vbUWcSVZTnk
RKlo+W8UWE+AFejHay2s+ZcQOC/gxa/9Er4dIplYO3EGUgWt5STzjVffrGYf4pqA2e45eGSOF9i7
84w2XvdDT4KzWql5/2XDvj8mjxtK7HoOR1SkdoTQ3qZ99uBAcywIU07Vwztj/i91nyEVQVcDroKN
0EkisWI1LykFGjQHdwKwI4/GbID5YxW0mYASVttSD5Fj5vZLcIgkeGV6aAsVx7+WZSZ3mji3Ib0b
q1N8k1pgSGSvme/E1objaNYLDJVUZW/5iPb03APnkw7Q5v3EwLFovSJuGJxwfUDKJfvyREybRb7l
RophL6Q2BlGQf45bOSUvkPVSW8SYfGWgz4Suzr+XTuWw3/yanEUcBdEX73mSh7AOsJWHwMK/WkZU
9THUdHEToK02w/PNhPqfTF6yuaeIhlczYXIgH3ZAFv46FAroaExwmpninCWg7I9uX2wvXQIKzG03
r6uMWftjXqgeuzRoXxosJhFHVBSC1wovX7lzbogfmn5d34fodc7OVydVEVpOUiUy/p12ZHsYJy8N
/ufwXt9Fpfov9FrLyhLpwWpJFlzfdSHWH7MLFRMoeJYdwKypMdHxCFWBwz/it9qemnJqn05D/DTo
CbATUYSV2SEC8WR7k1c/Ae6MIWPSg903JUqVrATDQ0TrFJ016rGxLd9/DEi+O43wEjHwKJRsYBJL
Wg2Z7SJ8okYPyKOvWPzHn8SAtbkCWZxHnUThwPev6AZX/s55VNqJ/qvfaE8eAStbdkS/Lo/KUtFO
TKS52NTAnvyaJsgY6ZsajeGkrk053kdOSlg6DL+CXFUYAh+R4WWh0KGswVPuC6RVY5eaBwu5E1o7
kSJNPvrjbw8JZ+FyfzSLxXwolQIpyBIsiZwq/P04UbaKcnfoCGs+pgdHz/dbNjrNUH2ng4V5rFw9
YKm5QlVsxS7TW4F8AElY7IYFQanebXNeEeLIY9ZPUa2Ib5ydD9VNH8yxt0+Hy4bFBHg8GEtVHacH
yki8z/r4iWHoFCDPdo8Dn+94Dp+zIPXZeXJM4jegoUE4gH/eThXnGKb73XB3sDxUVUJL/vmwrAoP
20QluK4RTZ29VhgJVEytJK0viLqFKhcG/J0BPdIJbTWaahRhJqRA52W+Zk/six5oczpv7O+v9oUO
njALEGdgb2nOIJgoO05h4kL7kSTNesMCE+5fh8GqUbGL5IYMkjN71au1/gxzogVcoe//wBxcm9H7
udKKJgQYPuGSWzWnlKyTPUGwVhlHKvjyAbsutmxpkvYZK4+p0JvljYpSNmoSem2QfbMEW3/JvMfE
fszbvPYxu+VSSDRIMGWCTKPJVE748E9AfiDQ9zKvuOgVAouKzY+9y5cFBDdgQQxhWBoCK8BAZmpf
OWA8eT+f71JDuGeAf41KZb8xx0Nli86Vmc7RXBkLUqYUV9YFXvBss6+qzuDMnjaS/4RHgnBSvRcI
2Sx6yIAx5wcuhgwmzSTA6SnsdCdPRhKpHiJWdoVaMprAG36/SWWvd+a31CsNT99mf0CHUaRDdKlU
nc9GNbhj7DYn0qgwda9OFIuL/zQvoeF7LS7h+A+gHGZ3JIyTQM7nybVdpUjk5s57I6mtjjHiFYxM
gWfwb0so4QhQdv+Td8rNDHqi178qp6vCPFb/JcscBB1KAG8G9Bcz6tacC6PLEDgNnxY5TESblGmN
sDT3X/nQoh9V+9FoEbi0vyFg6ApMQejGm04jvGrRsIsSy+UvRgDNPE1Vnf0Fmgr33nZiuVKy7syp
bWIVmaaKtXdYEbmxwNkutANpDKxhm21VIDyX/nXe5hB3eTCbjn97LayHxGRL4nDdgFuWonQd5Dy0
5McGqrgtEA/WP3tenSdfF6i8610mDRACFLs87gCjxVM2UqsIu3y9BWYgzCx/ylj+DnuYsg37PpB0
Pbk2+9StYOT/qBbOKeVF/mmBzWFXu5gcS1D+y8GG3XM2I+ee4xh2+e5E1aq6ca2rsa6ZdCYllq1Z
6okybIBhmvFPhJUY6BEilgc4GKNE6L305JNQRCBDi5NMR8yoD20tqetmICJt81a9jldwfswpOdYz
YMO6lrciDnwUG0xu4nYYGk8uXAx+sLclRCYMwKPT60Pt4u7tFAibwPT18yHknafDjEAu14/fyhuq
u/089ZilpVp8MknLVZXcuUziPsv8oZ08XcwbbBLXX+D9JBfX5LAIgBc3z3knIueqVjjhsh5vQ5X7
deVkKbbyX9nzM8AZjY4TileqH6GWmvDTskC+/5Z/tw3O0qlkDIJEvVaID3Aof+Gx1/XmxI3yab3X
WaBkkEDTCAqTe2UR+IsJkRHt2PttPfqi2zVisvViQxszH5T1ndlnoi6ot1ZG05ZFzGqPhmsjv/Pw
w1v9S1i+xUtzBJr5tVjPWqqw30eQJkYhHvywAxLSeQigwP5kolIjvD2BN1+viyyY7KZOv62h/Jrg
HMTPSN8yJaQvJpMvoCRVzQSu4Dbt5NcXAGyo70f+9SArBi7K852eiwwWRglHE4QBke2v7QNYOjZQ
S9f+pkjyrst4Pe+KMrW7wz/tDrFQ9Z1dJyuHpawqqWiKnZr14lVP3PlPW9JGT4+kzqFKeEUP0tQr
AJE0ltNj/GF/StX5Vfsugw8ue5EPf1+5U7lDrcC8J1nyZ8NcZ30mKI6LN8l0O2wIyq0i4Gm1/wIG
+gpXNOkNpSoEGN/mS/5VFlhg3TBLEW7tMD1BeQRWDnWlp3H5J/o8vBh7ExCu/JAPhCvihovVwaZf
P4ZqZnes20pAwFbFb4U9PDl4DR+zhogC5q+WuMLRdzg43xV17cSZ87I/PaBXKh/T10Emy6zKocJf
NAQvkbG6486G3tn9vLcGbQuxc8MaHc43lHrHYx6aDvAk44yOK2JRkgIxIqxIj2rUZTDWaF5OME0c
ii+GgKr2FbdrNkejVs3DmjH8T3LjUFhQfhlWxzfEn3wxq5PhE+WJbbGQ1fc17Kmc4nCRU50lZqex
Nl5QzF4zXj5gfy3yIW5t8D9l46Q1aVHCAgCQxmfVZMtfbdCD2cx8JdIZeJ/KXtN1b56kq7QlT5KV
yPeFDX7yyPrLQpB+qCxaEpVVwQ20Oa556XAZqZOONkx/F+YESdGuNzqImcVKO92g63vuDfj96jAk
TZCtEAtsoBx29SMuASEsh/Zv+SCnQDTU8sPACVyV5Ew0B8oS9FPMX7AMlsAa1s2Fgvzl6L7Hlex8
qTB49KX92mw9LgIRc7fT6YQlNVIcITBMbjJ9yT6Rg5esD3kj4JDiHVT+6rkPDrJRnGthRlKEz9ro
FiDmJ1JhzY2N4y5zBss+l+M+86Q6iXrIZpvUdf5qIGKZmKrXC75A3Hdy6f5QuDzfhgjKcc1KkRRE
L8Wssh7KMsw/pV0T1FatytnfUjgxMLVzsJCq8Rh3wEGDOswnAfA63bhx4cGkGBFlixppAYIPF4Yr
N36g07YkWsAgUmgeih7u/jH1BAH+NSNqTxFLBcmyRTmsYRMytdcTiMlHuQAs9uT5w7cfEQmjpk+0
vYqNp6zjqLhTU971AuwE+MEJyhbCS+zWFZywYjiNSffsoVZhjC7JsD4TAtafU7UpZXFsnpUmtKW0
2mWL30VtuwuycaNQtRtUQDRx9DJufE2Fk61ef3Ol5yp5gPhbEen29HLrCVCpScFT7V7Gdk7afX3p
oNFUAFV5Xm78DUYrhVs8DSYK88Hz6WQpNiXnE81rjgu7mWxT75yfd5QnoPPUGCY9MkbcHrC+7oj9
w2Ag4XP8/KkAlnL4hNeVYv+L1J8ry9tAf4fWj/L/Z3g2UEvya+29f5NhLUjONeyHpcbaPYdKjABG
HvLi+/G97RO49KvyI4ffm3+Aado+eoHup6L6+cCzpwsK/mxuZEzldm3VCURNAnJ2bGcBDPrvivg0
1lxckSROi+2qsGePRXA8wUtH1yFIeg7qPSWZd90xn9YkU9F0FNlzALf6nSsI8HAYv77pXP2JBRC9
2KP6Zg3ZSqgYruS/xbbXza1J7J5udVObBuECNByAi2KfRd2QnMVrAXN7+btdl6HiKq8Eq6tBRKPZ
LOuptJ8cL1A3+Wrj5N835zp86LmC8hz4ppzazXPNl0TbFGNX68JCQOxIuBCKdQayGOdA7V7MrP5E
HapzAYZ4nNz2hcXtvASDMpd/3qvMEw5y7umjrK6dNzcUsjDV1u8K1f0e19+y+3blnAIDxkfENjWx
ZOhDWYH7OpZgKYQp4xOf9AbSO2n1Yk4VVBMDCgaikQrK0d6svEnGn3wLICUGe0nAQPbaD0ATjfBI
K6obXLyRZ4XQs2a48WOXQUWdj9GKMYhl3mU7KR7D9x4YxaSyLzEpjQZOhHz+YqxnLMUU8bxaUWNb
JZe8deD1+b++n9OsBlICyIt1WCc9SM6zk+azfAxtyAsucaAl8ynkjTcU4zE6jZoUFXJX2o5pM8ZA
FeNRQou6d+gCJlcFEKfmCxZ+EoSCSzJZzbfiFpx3FN3v6/2Rx5ucUd9Nl+flsnoMjxcBIDznzIPs
tDr9USohyABciTJUCVkQvZW3B854TosUa7z10YBs4/ggvYTPA06IXhfUQyX//96t9tQxQ/6JaHz1
YVoEVoPb/E5A64L3dKMmzpnL7+fGTwKX8gZe9hi/dnBwReFxZusfWb+dxC8liRwH8ia1o2TxcCCB
Ug77uiJfd3D9lqSlvsJHBIwsE/6WN1e5YdvhnkKtNr7lqKRqdb6ca74O1fVelWF+CE5pw5Xi6LUA
t2/3ifaGgn3YSL79aINxOlauPETaO0XbFMIFjAbvCtlX1iehNMkCsSJYMqcl5Z/FU3wUUJXlUvT/
IoqkcjfMsC9aga0M4CDlYoaIlfjT0HIR81YBw0Cd9ldl5S1Fm6X4kHBQ1cWYT/g//WddKiIYTXUN
bkdO7S3m5behVwIdJnScibPCufqgkWtqtiSvU6DkgJemtVzElV6z2I6fPiWkAB3ZuZMsd7IKEOYV
L3rs4cV3qOXaQaC4/F8FNMJ6fGn8JsRX4bB84IqACYtHo26YU8M5LEyrWrt0T61kq9bo6G41+xrs
NEzUKGNMsYDqmBYYV6sr2b17bKBboU+70+ikeMkpaPXV+1CDEenCX+TZOrhc4kx06XJsKTiHZ+um
H24Dnky0Fk/7rOuag9JcGDqGD9gAUXbmEDJTk085vN9BDDR5fb0obubXCMwDmd6t6SVe6T/u9nmO
Dp5L1pC5gK7ulszbtnEOAXLUhbm5dTaxUA+mmcc6bHMyLEZtnlwHJ4r0NhcggWHEaC5n2RQduoxc
99AaNyJhuWMmN6J7xEv0dWob6Tmvx8wkaR+axNgox2p1Edtw9DK8sgVa1KgCX4cRhWnRC4KMtXhG
fLMf+S/gSBSs+QgM9FGcPo1WWwNtquCGufiGgxFZGD1Dh1/j2aZ7TKfMcDESvWq3Wxz9JeUP2LAb
bUrKrQi2FwSWm2umukpI3VMDgeXPjnneb4HP5m+j+Ovf10AOSlvJeHkbOb8i/kC4p/U/5HYuyfZi
q/PhIOfrmPMMw5H/LJPQQFtAciug13pnzMQmH94ZIm/I9/VwU4VCjF671CMpyIwfxYCc+8f1ts3X
mkOzVZIUTpeCvQXE+JO9cE1LnDuhTX/Nt/NbnjRJJfvGsVuUn8LouD8IYQmRZjIPh9zLKd+sZ9dq
bvof3SzDgf0AILXLqAt6TtX/eiGkFhw7gkn0HBtyGTmbhCPH2n6Gg1UrjZI8IiX/iJH4Kr/SZrr+
/ECElefVDZZONSV3tvPUO+RKrY/q5PXa9fKQ7Ffx3eXGbVLy9POKFEq8UI5LPSsZ5trso0sQmE3Q
bkgZUjEFWF3zEB6yq5bY7NmQQ5fL72PIW8jVG/fyF1NVL8K7jL8LrgowNGtZodILArvT+bN/475Y
VBC4Okr+5BJ67+1WZQd7Tx+H8KXwTw4rtx66G5Ko945hA0pNeHtQcc2iwpkfEcCCbIMZ9RUBtV4G
FYIwaySKQxfOHGZveRcLqfN4ixlnaxusBO0aYAQlqQubdBJkr1BjoKikStUhk8zEjPwp1nPqqN0c
9s/zjh9v3RkrJaBFAfphntoOxNaQiYLGqvAGnhv1nr2g8KVJ3atL2mcCHiAZ+YzMJ47fowfKd7mp
YnJN2Q/7fERc+/0hvfX6XRisf1M/YwRskX6FRdICV9O5aeO6MtBV26TsbYvNGlCjBixxdDsCEhZX
0srxeuHDJfv58wdG7ciTuvU3tPR2EvCqGV7w+98xQ+r63Kip5vWC2/eBHwD3upvMjx3svUPwLCTK
V2zEvGmBMvMHbhQ6ln+/Noq54tHbL4RNT8WVZQ9EFVK/+hL+00r6C2OzurSAZ11VWl0G5cMsbZXN
HhbMMyY3wRyPNvrNL2CUhA255WHEZlsrqG/ikvQmtLUA+0czE9Nuzbb0IofPcQfPFZSFACMiAGw1
IRisz6gLfzTmS8OxbQRKxESIGFIOKtY6+6wVEy84ksnZJqNmY/tXTvQ6az0+lEJBZ+5Lqx31ZfwH
azZMehfQCQJfksJaAWcww06IyltIcW2dakyNrIPdo+MlRjL0gV/b/vQ4ua3mzHWWLgtOjcsEv44+
UcNiNmvhRxd872xdnaiYbl0ARcwVcfdcZZjub1P/G1eQ7F4g0wcNvaZ8ePLvAyDX69RpSoqJ3UOc
8EZCQjXyezP/nOltnBcLak3MBSIxCp3DxmuC4/b6+oCGt4HICrZepeYyvPhogb0gl0Tb9+In/jDs
89DEaOgwF898WQMFw2Z3LJPIB8GRrARTZpT85maCuog+JtZG6gAXYKuYKVpDixm2sHwryIXvEHrG
+6H5+SmvJubgFU6iaRtniZ5GPYPWpnj3esWUplsHjjaBQa4qDgly3AkSGTGN2PkX2gnaYlUjKX0h
BG4XtVazbD5k4lUWo56CUO0XmHEHxEhMjYNZmJxq/hi9nn4DhOwQ8Xjo4Z9/6SGJgB3kh3v+6f+A
HC9Jk1HzNVjzb22soS+K0FM9undOgijpR9vLMiRbkPTgePggw4UAdPLhebsNfIOXXR/1dl20N6c2
AWuR7BkaW/Bq4x17qy8R3lFkWxdHWcaZb+eEdrnQAcOHIC4gWDDuJ+4mMeRAOR6G5ui416y94Myd
lxGhdgf5pSWE0g2wjrcvf5MeUPBzbtAgGE7U7mw2HozjTUELycPm3Uz7+gTLCTi/L+tW31TUhdVM
RicPaosQnpnBa+zEFofLyi+KRQojeLLauwC/sTU/Y7m3HjaD2j49Ttb8xADfEz2l+5xPJ+uSP91F
moT+Rix/E+3fFKZ2paCSbttqNz6Y9fzlKjJBLF6ulD9ghGHlF1OzZ1cj25Wu86QoVm0BMhcRgz0P
VSnBgpE2Q1StArRzERwn6tb0ZAz8Egq6ltu0o2pmE470VtY0YTMLqEGcqh5kb4NmxcnjKSaRqwv+
4UMTqfypQKgnGACHO3Ar4+FQnmJeXUAyGN1JMFbyXOFwG62dqDF7lvDc+sFyv6DCwPYst/iWKi1G
kGSi375tpUCH7r4t1Cza4cwrLExATKvzmTI5MH4QVXiN+NyE491hHf4rolqvMC5xDEGwTqGK7X+u
RTiNFP+ZVwtTECBcLZGbVM9Y6j4v06pE4KQdjvlMw8IMTpbjg/ij8N3d066y4w986sYYvsumoVsP
jYDPrbeTao9g4FblAHxmbennHH+cAfNOL5BymVaW0/vZEMY0HOHKcT8casn7Arf6nm3cvb6lsoed
ygX9Dn2A12GnpWcJ0TEw2+xiJoFqqtZzVpasdwDZDJ4OimZucOf8Pdn3AY1Is2UWP2g/+YqWfXUc
oyw8OYkEcL3qp+cHoVfUoGaUT7ILDQzLLsZ+ZOqAnVq+lLTOjJDDllrIc2T3v+oR9SfYDI0waN8o
4sr8pC92VS4Se70x+DmKVHkRJETj2GUqCLjVxGw0WQezdiUYKu641XB81EVoCYm/r3mBq2pKyNVx
Qc/rTz7B8DLGuAAY30txFI+khREeLKxz1Zi0U1bVJntm+JyeYkxGREo1MxxiSIRqJO44vky52LXh
+kxIiBMN4Ydk82QCpkHqIG20+6hJS7Pnr2DtmsI6ofpu/PTgd1D1mVevleeLXMJ7vFUelpp1DYKp
8WxJIvxOrWzT4F/MDQ7nsjSLeijTFpyJTITYCWayQYYK4yhVj4+l0j+FmYSAvKS7A2FDRhZQHh0N
q1Ywl3et1Exd6BJ0Y66d8vVdmLjVh9k5DD3Y1ADonG3QVJspw4T5WtrZED5puhVCZsIhXURKnRDW
iegKAblheVbIH90newkMAd7MDFPqBbg+nmtT1CrlSNB6QJ+C2rH+HurgjsdgOmeQUGVQoxI37n9P
Y+U2BNcg1eVsLfqKnPRrSjL1R6lvr3VGSxHAc+FHbzTx0JnLhG6r0ZgFrJLur+AU3kHwVWAVjt3t
uPklFZJ6b2NtH3L/eyEybZDgyX0Gx9q6KxXSGn/bm3vYcdLkF0U0vy3RJSDTmBo/AyTbN64337S7
TiffhPkPasA0JKbbOfZAPLKwo2KLcnPm4zimATMTR7U//wROYWm3osfRj0KtM9o21wEAieVsbQD1
QDvVLPYBA2IPoh0wPkKvNHRYZHZY3oreOygtFBX+t/9GqFFeI//MCeYqJh5mPnAEjHOndGcWMvo/
OA1cydQmpPpXmrxpLH/oC4TrJJ+VR0yh3DRCKIzb+VQrmPjYE4ZVyyLgsE7avKPOBlx5dDZH5mw7
pd9YwD+lFDyEI4kdZZNrY9Gxqb3z81elUWq5hVZm90j2f4nMbx/ozo8UA4uFsCKDoawFNFGp39hv
B76+VYDLIsZfx8w3S3aQDJ9RQKaB2p818iW/RgqeXWIiw4DMg4ExLFwUKZ77flSMR+RnbMoMgVdx
Or5Jm994MYmMg0PriFTMPKtRI4qVipJqbbjDRpC38ey2wa95Plxx9rWfC032A4hhKqqppBNhVjMH
kt+z+zjmUGcx3x5izDEvA5uPZVO3oqb4WCawdDFAmjoFQ0G7ue18cLUjd5I218DLPrBG3msMGgmD
ZGGbainwVN2/mS198oICBDkBQhbpncULBwW3EIfeuuxVCj0JM96Cu5/PQpA9ZGXnCL2bzmT/nHs3
/Bs4eLGJEusmmNGOSMVpwBDaWmQ48wwo86g5bY0gsl65tL1UPkQIjQtk7P2I++mqTL3xoPPsgkhL
jf4045xB23N+Fn7xccZzeXLf6IE/Y9SG9njSGkYSVXsBEoObsCVG1zZGxYKdiEigk7ERsNHCgUtF
kYdHVBSnmFYJDUWi2jylttVmdLC+zUNDEpvzA8EjHqhwSWEEeGOk1+xj58B8NgC/7atisHRfI0Is
uBDQo1mw6MmYXFwypCmHcW1C619JNcUhecSy2+nrfNc/IA8+oPNFv+5xZdECX31OQYo2tO5EmTkW
VsUnmjaXUzeo5+rAETBkebCA7lnHdQfyQHvf0Vow52Gd9eBm5xcEKerNutsrPXIALy0Z6UpHkrw3
mVwNgxlDIgIkSOOFh4kLNtFv5RiKFDEdNXkK9W1vaxIp/JsRM1N9RDcUc5bMSfBg6ypqSB2YFuAS
F4o+DQTg/hkg94FSfUB7whvq/BYSyDTOHL2BYSR7+H5RFFJ9XJGvof86SnnSMqCrKf3lCEIFqfwS
C6BSzTYrhq/1jmhNknpk+H82JfYNaIwSDN+1YUNKjBHHzx87Zj3lF2tct50/C8njl5Kv/dwY1JKd
QeFFWEy1KjOSCCYCRJxqXZNq8L0D111tSHbLpoF85L1BA+lKV+NhffVZXD8GcjSMuWPyyPuChjsp
dJS3+4SfWAqOYnmISB5Bewd+85jxYdy2LzdpZgDxtWt6K/R7wX5XpSsBpNwf/QF6ihR22dChf+jV
apBsGyZcQOsJuj17GDrkCelLKXVHES8I05ev2ba1inDlQ6MYoHvsAi8qFDIoMVbUD7hNw2/oPY53
NTbswdEYcWduIbCATxquZu6/0uxz+PuAYL2+m/qGrq4izK6P/bPXHDsRH1fUbgWPE9nMEWgJuRMd
xspT3y6n8l0si8L5JY+bFdPRNi62m+0x0XJrRwuAeKbhOla9/4OVPqh4TP6xjcmIuXW+hcHjG65G
ED8dM6OdXPkanES6KpNrZry/I81qzmehlrKDpWNuOK+74E9T5NvhDsFUhR30qaU1+3ReApbcjKBI
sdIRqZKuphRWHpcOb4uV+lEygnw5ASIY1AvL50zSsWgyiKOwdWMMcsxU5tU82n2ZwyaIzCRo0vxH
Yi8qCzQoONWXhGxR3K3lI+PTEWnRfKSDusd6Dkdte4ERuP5VpsmzVBYxbPTN+6FT9Di2o0kXzEVJ
EzRFpqP2xAvyMmqF7ahK1+A8ZnzNiI8FcMTgFzMF/FQU/ggsCO28l3lap9/y3iiz3KWIiPUfPczk
VLCosImavZpku+8ukH6TBlj5gUCxYwSNDgXgq0klwW/VzuonYlV9UaVZtlxbm+BV+MD5rHzvWJmy
XMsiwS/HeXMibcVTp2tIiTdkQ8gm3APD3xKghHs1uLdtCZXnlLR3bT7ghKl3tkJwtnv75GSWrhT1
4MSRa0Z+8x8ourWV6qShFon7Feqkmj+XGapvxefCvYXZGOZGHqwaLKN7K1YC8goy19hWx4rpve5j
vWo15pnkq383yQUzsHUCUD+SRKNUfvJy0u3NfmGybHEEkpK4x+v1kuRiIlHFIY+R8/m2zn2xDAV+
SqtZ36sGUAMcIPzuk9OLi25wKcTC+rPqeDKlIWzPcPKcdaA/yXr+xjO6WzuNEny7VXrjZ5qrvlGB
wk+LSyddrJuMW5998+Vhh2+wYqNLaDzX1vcNp1/JR7hc/iCcyOi/VKXRFrqhl4QOFUOxyzMzg4aH
CGQu1FKVXk5VaqBhDyQxLsQJc079FSB6RLomtfsSi7H6Knru6+ldG72vIbZ9HWuFO/f3m+vLPFLH
fmzqudDSub4ub4vPUqJziM/ZkRlxYVOesxtIBtvjbdG9kb3Ja5c7thaAHc6jSAW52ig+0mzaG16+
n7wKe+9/sK3rZzOACYMVpVHIs1vtZvjxZyg0jJRkquwUexyv/JNoCnxabq8joggT88ff1vvNNHdG
nTAFbT3Zz5gJ0umsFDzjVAFJ9X8AtKys3JLhBbdQRTxVW3bKuIbiZSJ3pqE5bKWvHcYUPysGWk0F
XRAZS8j7DinZ9WPmPI7CHWK4y5USoi0XUJxrHAoxVmXraAs7Iq7F1fis/AyBKwyTQ8Xb+1mVzb1F
PDKK1VNrpDILCFzjeqUgXog76hHS8byJLbl9cw7C6+zBnK8tSKFzNiP6i57plMYthrvRm65LrpmU
9FzAPFgx9Sd/pUiRX0cfKua7DQP/nZhVZY5Hi9mRUabXqmXtVcwEwabRlfAAybaHhfDqeWul2746
ecX0qW2Iu5kip/GoUhWsgvTENqt449gjOar2EqH9EvEhtPI98fZIcsFe5eE8Dbx2iMF4AJIdnxcY
FKwq2pQsJ9SRiYL0cnovRszQOjrnofgvZQ7lZleA04mEARMawSS1f8feRpurtlq01Hkgj3vdXuYc
NrRt400uLSjoPn+ElPqT1RqVb/vtaipUDls0XayRJw6TUJplIbFI8FfYdc+IA8K1cRmjbpbG0Gjr
poktvaWGWhD1oqVMmF8FLa2pnf6ad+x3NuRn4x2XqcxW7aYPPliMf8zsbAT3owCcBkAMu5kjs+Ax
E7vcsLyVpzcy/c5JAGyLm48t8qS60GBkrSWT2JskX1nqjEOoCfSvwauxKwGIKEQ+b66QzIAzvUcU
5os52l9FOoHM0aw2IGxKuEq/AeaWNgcAfxbNdMLdnorEgzCovJ/Uh+xqsBzDsTug4K00rVUZpscY
GJMfFqmZsXwVG7AMicDVw2wEynpQQaNngv0E0sPDME9M6AolO3UHYurUrfPs7SYmt+uSVN6YTfO9
XQwo2FRLa6MW8N3JLYCwRESNVAD6kkx2sHteb12VWSrj2L8/3dA3ryqGPUXAzslcBCVNrYoIq0FR
eNQTRHzYVH5cO31Ts25OjYHnMiV0ukfKZXulbe6MlbFEMF6c/Jb1bK92J/0+UGB8VJ3Xw+Ed9lZR
x3FhYlbLGyfopLt1GtEKPZg6afQhFVmf+eqT+fkRQqGPs3Di7aeOd7gTes+bURFa9Dp2x9yAuFPk
yW0AyUSXr70DS90cXqcJcCM4fDptrjC8C+imIECEQA3ayUVUULaPK3z4yWHG7x5NlrkX+YLFbVtF
D2Y5W1CWF3qJ7edSMqfJyameaE7MieAwhj6iV5AKbxK+9Wp3/HTy2AATOXMhVvZ3oG5vxa3X1aIx
dSXoEpHkRvtpARcZI38EXFckNvUCjPINWT+WNYyHYrRxWsXk1Lmr4Zw6cC2knZDmsdpRwyHVBNLW
3+fKFg3p0E/fUFaim4QpUFyZEQGcGVzYTKc+XX+D8VwYzqFqrGoqjJpC7Mevd7fSkLM+aYIqqMeY
BFKukaQHQKqjOags36rOR5rAHLdMZukA7jCLjNU/4VKezPkxwW6OOU5gcmDiz7TFLCzKnm695Vhn
4jRO+I2J9/T55uUDsHuxtUA0FYmw2DyjBaqrbq3RX2QpX5lRNTxESoHG7433SUIWGd1RNH51mYq4
wkJFT/FRBq8w/MNMVAhG7F6cot9BIPjFd0pQ7zFt/AwOGSQXL2h3VN36d00AFCvXIq7P7h+UOwNd
+RBZ9pRrUaGHPilhs3iPKcX8TnUAmqRExz5sdnul2rN0B+J6t3cFCg54gCb6WdnRlqkojpbvHAyP
KghHgSzDpn9MHW+7L0O1hQZhFMc3or/bByCNvv2M/ykAikJjmpPgN4u9rK7fA2eL4RCvW8JgauDv
/N9ai5Vp33M9NIkETI393oaUkaEkh4XR+iQTRza+/sImdOaZ//h9hmVHNwfylFuKZ3EHuFF/eQEh
e6J35ZXKhldLOino38/tUo+KhiinAQUzItCKcgSFk/5c4t8mwo/rB8lDA+7i0B/x1gQneqZqGBW3
U7zJLWb0xpZhWGIJD+0bbgdcc6Co7hskP09qy8Blmyawu7fc+96Y9P2GtD+ulI+gpw+jsY+ouozT
no7gdnjFAGepQgcTusRDi+MMZhYUqOaNRZKF69fBDmODWWQ3OVpOkjZuxXnB+gzhiyJs9orC7Gbq
nwDtlS+qpRR2V/TyVLnyx3zejzl/Ma3Sj8Cl7WDptdqB5QFwMTijJI6CPsjb1GQgERjtDljeR1/7
xzIteYjh7k9fO21vOh36bpPMCqjLIUdaofVaNCHUwA9wyRBSZ2x4IXXWtyWbqgl77+3tr/TJuX+/
ukcrfqtcMVHnAVfUJsEtNYs9KqgcmfJzc6pE/ynZGJ3UeArIUD+BWUsAJXquRmq0ny7yenVg6f+0
R+Ra5HBcCPWwDlL6acidkui0ekrCWgDSAcJHIfEuCHEgzWfrL8U/+OXBz1nphg+nbUdi6qyp9HaA
E+vM6JgcjWlmCZW61gFcp8dGdbJyo6vCsm/x1tY3OYpX6yJZlP8SUuNsif0UP+WXwEXJkf774s9d
VVSei5S5vnrXc93NidWhkNY1PLGuPJR3C7acv1A+7wtxzL3LRUVq7jPAGNhgC62jCaYwPzEfDWZr
Er9CKY5W5A+Z9iR32mwJlVh+qbZaBdqYIhT8CFaxvp/nq/vs+uc5GlzoixVz5im3XHdPNjtqko+w
ysYjJuXfxfOyXKckAk0k0umfjf15KZM1KRT2dys/+DRuB+O+ETHfi42RaE1C/OQ88zWs9/+g32B6
8yc+HboMlwcg4Pax766+dimLe7UVvPThTQvDfUwCWh+l0SkqNnepFfsdEiOaM+jLtmWIu/3w1rRt
ZaPf7XEBzO7c3qwefGvgy7HTYUesuN/NMSg6YdJkj/NXYpql9lPxuKcq92MYtWFpJGryzvt2hW3J
nxEzaWxJoEo09iNpBI7l71Lgi5c61kSX7ApTDR8G31LradahE4inrUMhdtk92z2Or3Wv3smEEtbw
msaC7ycN+5yQuNLE3JU9zNb3nkYAbVcTzSj6K9eu22qoTy+d3he5SJ5WZZM2VgmjorgXdTDbxM7a
wV0jvIciUKfks6i2MLzsjNQTpJ5ALijGIARktiz/iVYHr40n8RfsFYD3ZdNApXTaeYccL2iCWqPV
6/qHwqr1uxDVr74rM1ZmYAuMeHZ2xJlfprQZrQ0vbwuwsaIuOLYx7Bol+v6D1qauGsTTEk43uD3Q
DtITiPrFlqbYWoXToWkk2J2mmfLp3Q524+11nxt4qM9TCfzZyMuIN0o6p1isyLzVny/thDD7j7Tp
7RGLDoJeHOAIYD/hnAtDlRQwNZ6I/aHMIAAbvsefXdMtde4XwdfBFq35cURK9r2eDbvhI8+Piaee
t67wZHxiMfcdFLH6oE1uYXTzimdioDtjCqjNPqI4JJOPwwbQrJUwTay2K32r72eBidNbBTEkAFKd
9DkssLeJsnCaV28TwJ2fIb03xtd+pSwUKdYV6Hzgc5kQ+h5npPz9wpnWSpAGGjZ/rGT3mVnEcRVe
KCxBqdQK9BFVP0HXTJS1Cq85oWvFMlX7h86X90E+qsasU3ndBvTlGDsyny0uGFuQOYZ7+5K+8+Gg
er8QfSu8LHEGc2RFZXYKh6pKa2N5k4LCHWINxzEvxL5PoxVbl9cKm/Talk61fKdV8VB0/acDaelk
L5GcoyhTiEtDO0nIleI+5vbpHJcRtNnc2eYvo3x/ZeFfNGE03uN6CTTnch6VJaxSXSZ9QZcCFgV9
IoTShqkMZpQFtS+8QgqTPOaZbZ2kd2Uev9SFseOLwJofmgOkqJiAdFp4G/qnqybr99WXmWDVn3kL
tLr2AqeHzkFL/YolHcBIE6TVS98HbITg3k+SyBijJKED18rFQ5fuz6EloS3dzy7KWTGWZKo7/aIs
x2TM9ECiFWavvQSZHFs70oObO2T3hq+KM9dJ4IVtugVIkR0z78VyxR0nUbNUxJjG0CbqInp4pW9m
5fwLNhXQ1HqmdNOG+A8VvONeewrWbsuyLn7TEWLplREE3hOdSqIVhgzBbtAeb+tYFk3JFjfNytHb
Ap2IiKQoJ1/fjNyWRlX+9YiNTDztK+Jwo5R7TNN20yjeIm9QrnkG8zG//5LJwXmYIGD+3D5JcvQp
VXeu3fWkqCdupZcI8kAQXjWhlfUConR99HrQlIpIJ83sxGwRYv+h6xNtfmf6QQUQyEHLkEDHDPuN
yuand6FeeHkDcAFtK8UZnDBDP3NP/qXEHS4BlOsIVuL1U+ZNI4TWG9tVFkXczDj8A3douSOjMz4m
ri/C2Cdx0aaTvSiNKptZLiWOoiYR1ty1YQyzSSfyunbnvSgTb+cyveNdnB5zOkVragePjyeBVIXh
O3Tblx/mjrPb+eso+e0d8GL6y410TBMcNiNHtyPoBMnWqO62LqAYMGTpw8HWBc3+LkNIOZKhspBp
QCNQ6Sf3cEjQCB9K9k7wQVxPWaBrp+pa0h4yP3o1hWEgUz5rI8QmKD40gyVRDiORX5wINyfHCwp4
rCb3xmB24J8givf7dPjzxRytweCCuXjL4ROQBLZ9mUnSJIsJGZPuWqi6o8pKrEuD0E0Dzf334VWq
mdAOZ3lw8Tl02TOGugwRRxYhmx8yCcr2vSv7xoe84lwQUDDg0ucdhLjry+OOP4A+ttgMcw1cusaH
+6fh0JI/t9iuOM33OUdCABM1ZJHpsR0JqkZ3F1Jpti5KfdHHWbq4hnJO60k/JyXlxy5Oi8k4Fwd0
rhh9gW4ky2oljsjDQBH6q92A3gx7RVi7kmp6IRpoqARIRYuystLZddyBv5Ya2wEOSZtvNb+CEHIs
p336A2NHZjbhnux6Ft+/CR4m/13ZF1WM6ghUCWvf+v1Q8mOcoSj1+WRJilKb2CjDD3r06vgEAP/i
q9FPc5E8bco5IHYTWTJGq7TtzAjSgPYa1lfBwl8pVrC9nFS/RaVu0VHdPNtBN3oHQxk+6CIsFS0M
98XYiO6S0bFpLLVlLYhRTVfOIm1j6z6BkvmZJWj6V0sIMbWkwmD8nhR5xDCTNNf5kdOkrcHgONf4
jR3gr8L90O1hdHUhUtZ36zLD/kod2braNN17YXShVwuP5MNSBSqReWWBQQmUymnSppy6hCI6Y4GS
bsq77jyl/E2IOa65oT9N5kgF2EX5v98CKeLTI/sAs75+el9//gSyHtkWBN9hdWU7rxrmgoUnTraE
qYw2jLVnjUTEgKjnLx0V2oXtVRdrTBep1op3z4rfMHksUGO5+/2ozebB6o2BE8A2zaG5fV6f0DuA
r4UcZs3kuNu/YQJIkT29GkujBcEyC85FzQ5VSIbFTc5XbXD11d1qI9h+FMjJgW6WaDgSxQBQeLmW
8UCh+I0tjCmI8pjY1lJ05hihGNsZ9xHkuPxSLZTa7Fkel7VnwGkh5S23+r0+ssYvhR4V/f1Z47J7
IpM3lK+e4s0rS/zznylglzQbxtJNQ1rVxcwY/VWV6N7yihZfHr+tST+o22gI9oqaeAqYCddXMEVa
PKLrNZC/utNQx+HeWUIbvN6292iyCYd/sF5M8zmJcCw6ehVRbs4x/wBpqpP2BerlJCugLeZnR6ah
fuJCSTxB00zRA98s9nu/qz+w7KNOedp++om1sHRIv0056JSXX3Eq+75k2IyzoJf36pEegwTAlKmG
eu9qzHyGCx58Mls7t7zNzqXbTSBDTN7RZ0580ragpcW/V2F6u3efic7aB4hz0GQXrEnxADBi+dJ5
phs4WUXelJinuxuwnrC/S3jRbqR+zTmJ2sXq6ZX4faw9MHiH2yq02btYhvPFvN4ctB9NONZmwcdt
iNLnZjkOxqlCfGzahBME4s3Tud+eWUMFH3VFm1b/Plkgk0hKy1FxQ6lq/xpmP9L88yJPeQbX2AbW
KZMS9emc6GIfL/ePFrqubN15b/cq0ySQjeQxFJEgPY8fjYfdcdqcg9ctOeFAW2f8rHcpGbgJI+By
IlZfcbTKak6DyLnCiRs4BlAEs0iY0JckALTl+Nl353uZVTC/O6TrAqWfsV5yE4DR/m9mzA5d/xLl
moAB/dDFJI/I/uMvNSOmQjhkUVZhNp/X0PCvwTWaqrz+EqzqplIY0VDU5TwiNRRYobnEddC6FwlD
BFDToCNAciWzZrIa6k4qgWD3E/f2R+nMwAzSqZcJ0dpGAbH+EMETXbhwYfCSTf5rFi8fYwn2ZAUd
wyD5a8mYn8TaG7cfnvAODE1Pq/yGIsxMFqvHcWBjx+yFJcfQ1b4LRsQCrgSKOMUIUrTO3xXnQEg3
DsGap8g2jo6RQA71UUoCd42NtG893LwZlB9ZFLqq09gkzbP/l5JAOzVVILl+tByqytPOPyYslv1Y
+8HHwFE173feQMC9RXaAt9lnMxfr7x76H25HrBRd8zFke9DTZklez/Qjl2Yq+FsfqwQ2GT8zG4By
FMG2qxcKIykc6M6HAXhLcg3cPZdBnSu/YLh6XE/VTzbSVbrRol7zJS4URHNm+1VdnHO/FUxbJ1uK
kL5b0266TFlvjrTrZE00lqyDd8UZtKCc2ckaO+v5mjqJOOUeR60S2Wi5ArIQvCOx0iqd+LELDN+D
xWHJviafNGzY44wKoccCcB3tsAYwjkQtRrgagbhD+nSiwMPKXDtGGOZz4DCRp+p4XywyFXPEm/mw
d0BOpfqzbZIya6Os5oQ+di6RV6TBU57xg4JXeuLrIuU30rRYlasGA7uppZ3aggshTaHGtqW0i3+d
v7D4e6qt51XCTKI3h+L22A9laHWemzd0hPrmn52UPxHeCURwIZ4Kavm+Xe9RzprH3J01q1lgZFTL
Cox6kFek/fNJu9F4ckSwtjmldoErlfgCIyydlDIkc/3sqZIxZgcieTLz3kbtXUIC/PWrveDiGWyp
afDsqX2no+Jd7BBWn4j5kh4UOyMURV2mC3M+cXlG2LD230Ucksk2nk2jKBxqJfzjepr/pcxFqOgC
NABAXj2sGzKz05ftbxQ/tq4NTTSgWVnsawqcUdP/scW33juXY8+Ws9xhORItLxrxzOWEHzpFAuZI
m1+hzdI7htJjFyuz7fjiX0Hf+obu7zWvOdDPymSrEPhoXqSfS8LOjY5qYoPrmo6PctQCOCvZr7PV
AIsdOYPyxehhUdngJ7P+gt/CoaXFNtgkh/sH6YKw0QtdtG5zIP9IKB7C4i1IfNAdwmF+zJYDWC2D
oEd1Wb9HAqj5JTS5k0nLTgTOzhg9bIO1eNzNInGIeCKssZM+Nk5flY6S5IzOV8jqQZm96Scy3KEU
+cKeQ7ue+KH13JF1FCEdnPn8iyu82A/bQS2qRzHMIy3kcpO/G4uJQEZBsaQBiX4gzNiZQFnb+JjQ
JU4ZYeA8S2s1lhi1TKS//Z8ABu0R6RHaAgOOVFp8Ap8Eq6AG1V7izdbXzMcq9Vso32VtKFFRviQz
91tt7UGYnvGcAQcqPDt/6qjZmE9rRGfHbcKwNbYzhYojHd6cP3MeeCcAR/6Tm2Snvj+cCH1OS3XX
QlCLRaqmmcAUA7ktoAiSl4ojlx77HGPanNOhUrwTS3FqSecKa4Ixu5Y0dOxsUTJlwGbJjOK36+Dp
EdKv9JW1VT5+4+qQrDYkaMIuwGXEzoZnz1I0Z5WEQ9E0nue1vUCqO3/pqSoLAGm0uaFiab24ErY6
AXzjIgFQAGRWkdng5acHl6oaM210Xd92rgcwHuniGZ96UjN/A3OMS+Y0Q6ZkvXE5/qzrKw2ul21e
rUlHjRQS1zQm0HZw3ol6iE3ajRnsroYnnpx2sJ7cMBZYwVnVrvMQXlGMfTPIyZ5qn/T9Pk4NsAGf
l5nzYJMexDxwseVO05KDueOqoXLNjqGnRWgsZJIHTmI4UZycxPAKQt4j/2tdzMglePpyyRM2sNfv
FIvQWRUf+kJ9O4E4K9KnxWiy4L7DNyxNAsNmiIBDmwKQcKUuU4TVuXUesH89oH9WdGdHXUXLI564
uTG7SEKo04IoK7rvKaITDOMr0qAGaVQQdYxSAHNWTYOCEXCuR/Wtabpv6beTI/6maqQyjwn5wLGO
QtieItivxoBE2STXLsTFqk7qQgxNVoL9zzUfu/qrinW9Mukqfl68epfsbDTJDRb3Q4n6UPVMfNrJ
IVu/3ocR/T+8gNSu9bSyYpjtPYHz1EVOkB+1VClX1zd4kXcNjNLsoEZ4fziRjCeT4XuyxLmmzAlB
KIKjwFu725bzQ6HXtZJNHfWtf97RjOo+u4zFMUC/imhaGsyq5FZB9Ga2ORzeGydd/59bJr1ejgbw
OjxfV6iyQIW4ubhsAAI99wo9K20pwMqHr1oMPL/SqTrtI8bDjaqJiolM6ejpseXBs8rYIm0skhrD
NclhfzoK2MtEoTtMgwbX10S9E5ROZmYemBlFxjnN1gZiKcgor4hPgPYqGkLSVAH6D8KGvdgengSI
DHP0HuPEJ3F5ZubLRveAWbThXsLbpbOrreD4cVmX++bZqMVvI0Q2cTfin8yZlTuQybvDMwTJPcMO
8Zt58dct6/YuCK82Ekb2K14Uj4cgq60JF93pXifVJXMSUXzgPBboB1aq04eQADM9DHfA12kERT6m
XUsmno54/yhdvKLaovJ/r3qguqeBpnjHSHIPcY3up5tZs7CDDxIbuRfs016kOsSCrv4YlsYbS4BZ
f9chfB76IvpheT9DTSbOPlRugn8/o+S0XLfNGaShpGlnLz38+9o1vbXrjhMvcOk8fXwnLpC8qzNf
QIrfPRhWrRwmqy9c5HeIZNfdeTPj3MOAP8/hSWEA7AUVZAby3wQhCiZ9ORxyTwOaHamIkDBs6nxM
/xHEpHVEp+bABK4SaiYtsN8rkRW7dRqSp1HgbHjZ+ecas74HQfLNbILENuaZ9vcZjpZxCpNnLz0z
G75X22ETX7Fbe03FGpiD5QpuNJpKtP27Bv/9HgJ+xJEVrggmcSyk0eIFrkNDp008h4lWFnO6HF4O
q8kPAQgzWWjuDwTvI0/STtZHmD2KcY7M4xW47r97Qyo3892X+Bn5KBgFmrfI+BmySl6JEZcD8jHO
SbDJwxUJ450z8ClWI77luXtmPKO3hqwlqNKPgiRLjDsRWXJxxp12PlNtLbnzOJLHaMRaY/rmLwsw
QjPnFEFEs3HTcaqW+vLiQu18AWmw77SWgLHf+/UXMQfNO5c1rWPwUS3f8mH29/ZkTtiZpXV0Mbdv
qrg7+tGq09SRxRqj0QIaabmOQdhQll6EnVoCsuL6xthLkUzIuxJo0YahciksKLTRuGbIzyxQU+At
kVXmQ12vo+UU6J7GBKrhGWg2/r53HORyA32H5IAPowCi9M8wJLg5KoqmObPV2S3129UCG94W3AXb
Tm6uJCiUwAUBMK+JrAslaasFfBKbFbMRdqBuDh1OqY7ulF3A/kA/5QEYGEnWfhHCordpI+nMKM6f
Bc+S7Vlp9pLCJNuvpUptp/s+YaxSveR0DoDiZuK+ImWDJ/+th0I0zG+EF2hNeeRhodFM5Tn+O5yw
jK3T1vTfHbSEtX+alxaJsfPXKU8x4ZOC5J3eb7N6LdvFmyqv/xyFHU+2xkonR9w12IW+NJ5aa+mX
00WQrauQDGPywodSsSFCkJchVzgxvM0i6T7OK+WudrHCqPoJFz4sAWis7cwq9uH81uy1DFE+svDT
mjh7482mbBioo/uezsZ652b8a7xS7HYsojeGZxL2Jc9D9Z254RDIAozo0Tpzzcr3y2z9uMu2KihW
IY8DurJdzkmZ8ubxWEJ9Iv0do3nPpSd8bylvqPSHKaaUl5XrXeoCqkhVckF6NIbGp/jCR6oXZImr
e4FlxapzLNI5Qnbq6G6E/RJ86lI/xabk5Xg2yZLKS37WMBUdNbKOPS2PjpMIi/4irYEwcxVh6jIU
sYAQ27ad6k3vtoNNM0Ms5VXTERIjLG5cDeInIChC6KcP6i8b2ImOMALedwD3Rj9QH/e0sWtY+pJC
wVVEOVIk3a48L790d+7Gd8waMrHqL+3SJyru+acPM0FsAoaSeoZL+33NXFVFWrt1RHjetbahxzrY
dXX3iBcZ6c+UFxb/A+Bix6N9OznuyVw4albeMhjohE11PdcDrcEdcaabRtpNUZDUGbvm/z8D5C68
KGy7myWDz0tDpPOA6ttfTaiywBcsn0DGrksJkvzrwlUYD9q/Z9AfXFwc67eaHp38ABmL3IyvteMy
Vk9SBZIusljEQinCtDaz1/Gz67un25ti0lEx4QGStmFYB0baYc8uxNUPpzFdKoqsxQJNTx32E90H
sWhTdeW5UmQ2cvo7kqQnI+A4I2RpiIrwGrL4Wx5BXSmHLj9Q4Fxy/+lNhAEfZAFDNNcP0hCblOYS
TsoZdfzCH6XZQOz1euxj8944aOSXSiKYrUR4t5pUfJP9K2m3ddWUWCwL7ioPTQRa2mDiFF5EDgnD
tLwjaM9GP1zcOAa4H43kjQj23pqPbRkqv5W9Zlu1wxrw6G3sQiYwLiV7/IX6OMEeAlTFyToys3un
RKhL1YcbBpcJJhNl1aTAnhbvNVk65/L4NTm/cO7a9LbWwo/rz+mESP0HxaSr3CRL/W8EjiMOIJb9
4gl80mmevKQS5OSeBrlHhQIiWfR1WRn7J/Jg2BFXHTDTTBwl9Ih9d8307ldl6+ViAYi1XN+Rq9Cd
U25xAZBOI6yRgoonQWe8oJhWfmi9ui8YY+aYRVuoSTTONrSQvjl4IPjCJF12RNIiD8UGfrK47bNS
bGJiRyiGK7qQAJGlhSC+TW1Nw/n+rRk98gNBbC66fqOcri5tJcWpEvp6T3G9MT8FbaaoL8rhyXy+
n/Hr96QqJ6ZYLmKs4ISXFeRGvRMd4BZ1R8Kj40X3xPhNthsroT3Swt+NCW9qIx+FdRmiMWi4UM00
6wIduuPUZHdpZNfjH+bC3mVz0DYvLv65a6ur5BVZdttDsjXCDqGKANpJrTjko15MqFxypU23BHSt
NSfWduxo1nGDkHyblItRw/UQoDIZS6vTRtJEX7Bo5nmZEZqoeBH+OIQlsbt287xXdKk30p6WzEPT
yUMiN0otRBZ5ZmQWy3RLfLDfrxh/weYDeCjlO4g+BYNs08Okz+eXzesX8bVIjWHvEr43bj4cbM6Q
YFdyZDk6ge0HMPL5hHcGcESVcSjj+br9wb07AZorqKnBSAlWUHcwQOgYTENBEBtn4n0UcYfySKP4
Jb4o+NB06Js+ImNFolK6KTVyI6Dydhf41l3JIVq6ttwJ192Mf9QBlAWqYvjmotpr4NWl2cllGIOP
r2hQqBuzaSaPjuZgpIOw1yR0IrUnFbdCGVOZIFWpK7jxEomZzrjHp3jKr8TM6cgwmFpVG+d4wO/L
n8IP/08Y4Z+LghBEJtc1gJOVDb2uBkEJi6xVZD4uptMeYTb4RA/Tk++ygkgAoh0gCgfZxv4kfX5n
4Xb4O/1EZlJjvSV4e/mn94U1Eho3x4pu3p4hwTLPaLoUmR8VrDfbnOQGr3jnuQdWNhKnIiWpQcw1
hA8Px+t9sJCdOVLdk3qE5ET4qNyVccp7EE3xrsA6HhFvuTgI3/Gl9mrpYZbHGHsDkPP7cw2N7Uib
Hm5zko8FH7eL78vWGJQcG7KlaSeAvzwHvGjzZP69THseTa7tBtcFSP+Y1QI9d+K/mi7kclDWH5cL
enVFFHlR8isJsSYhEeQIO/tw14xvIzvqzYAT3iinYP0ClZtAOIWhXX0rwoK3fIecab6CQaVtPRVY
iLmEnYEG6l/sTZmaRmLyBIbiMchPuLPgKhbs1vHZmcJ8EfdiLKR/h/HU11qpwYRFBsjL7rveVEqX
bTDvc4nan8khVPIv6d7fbf9rf8vLPywluJ0pJgF3qlGmwTpIKOyGcZI6eqYyaai8hrWCLhKMJUC3
LNdVgVPXP8hfEHhO6peeIqe6VXAXm0y4HLyeSPKW36JdNhObCHO96xDE4qPnqcksRQLOoZxP1yOj
EWGqqHrpczCSoeiAxl9xKIaAXRh4KzruS4v/4II2iNT1DFDMv95VYIOZsuqlt1tJv9DXKhq6DgW0
yc5pgawQA/YMxdzh5NTA8b5GXszWTtiJc3dqqukJcy81aAxW7v3sh9fsX+fsgVrF71J9q8Fe0Ewd
/exaU5v/163M9hYfZfAMuPxz91vVY2gs2DnwHyz8Zz4mVsvC5ydrq0HQDhXclP0yUs7QLMpGbNEJ
yJKQ9qMdKA9+NLJEGZCzEz6xIP4Zhu/1NCXgxjJTjyh1B2hvEnRT2pu/HSaXSV1MfiQ7cmxsZQTJ
5cHHHmqV3nxbevX3rkpc6HvoxAXmq1D30IwgoHrS1R+4vF3q1Hkve4mvwhQ58iBb+15pfnF6UAgC
qm0PfEHHSq1xvQ5rFuWfkktLgTBIJWI70pviBs32HpVSqCU2AA9/JmZlgI+gtd89nPiuAAN3oTK/
hSigYTxiYL59kq6G8nW7U9BnIyK0uuesBHNLA9c9eKcUPB5nhFtpqsTQfPnCP5m+9cFQ9fiKhIcu
CEqaZ3LjD+Ay4nL8JLppdMhfhEq2Lw+QvdjC39CVgf99EzBeQbLjMLpLwZJ5BfgygB5zAItDPg64
JZIwj5Pjt1hrsrf4/W8vWw7cZc7zR1i58d/gYZlvOWZnHJZ/YsF5FhEDcwNivMRkmJDiW4jsK55t
mldLi0M83X6YSiHup1D+9EHi0GmLKfgTSHbSJTEGu4FGsCYt37EGXs19BiVDQPi7IyseyBjVTGEo
8Zqs+wKnXaoaLMYfvufiMgxQPR/LS9v4zuUTx8EyjQ2zMmXSy9JDJm7lEk34n+X6JKbIcZ2IahT5
HyyOQWOQtfz0smdbFmok05E+CH4M7qdVUgiYMFjfI1ktFwE1gdAZMgFpDAnBQfi25bRguMePN+Kg
AsUjoks/D8eFykX3OWqAc/vg2CiRFl1ktccfADxvliTH9Xbz711H6r0VJHndDOxA9DtBKHEy+tCK
3eEnwz085O8AsdRY4mMFCo/ssVmF7YNdf5dOUj82s7ibKlFQtIsSWXlcU/3ObgzY6AeySx3ao6Rg
AnnRQJQGifJdSAGBHt9tbTHLz/7RqhTL3/vD4lgOivfsu3MTH4wgYqG5qGjMrH+fCiAqkN1mLIhQ
qJw6ZZSOKSL1hpzAsii2PTPkFyyMTBJv/1zPjmbNpeVmTNuqNA+UyxCJKdvGSJkiAzcaubdHluKv
CIiUCeMiAH6gpPBtMaxNirdOF+VFZ4jRJPVIFTH/CxwrLtUV6+xE+ZoTMF0tQ+/ugqX2zEyow9BI
lceqZ4MIl8ytlcD+JzoteG+JwNwEOti79V9rqq5LOUIoesNwF5++UlX7UxGOz6zR2yAMzk725ebI
ka2XiS+Rq7fY6nFXOdzvidBWpYL7vBc8Uq104wPThsKpResv+6ifvB7gmLJTUsX/5rnSNEUit+Gn
jT1j+cMQagjqA1CYZK+Z0V6/IWD5ujXF0vXT3Z7Fa7Tek41/qwHWqWBT1FuT/JRmU2xuLz+5hPgE
eY55Ax5lsBYdNyMqDSbRymNucXPY02TahD/r2aHWmwnBeHE6/MgYqPsCowwcekK6Xp1sDGOCQQlg
JIFBXXCFO0GJ+SbP64GcT3+oskElVBMmNaNDt36uaixWl9DLMc1o20VVhTIyJip3FXPswKPeS6iT
b9/yjqyOHj+0juON/R6J8/AX80L2Xbd+Us/A77vTc4wxvtGybsWEKEgxxLJv6g13W8whNHzdDhHp
TOR03lsMHfUBeX5nXFg7o2CiCsLTFN7dAoHSAsR5t2Oh1oPkcPivnkUX0o/gGGHER5zpdy9P0HL4
172QI+k/XvblBebXGzyGllAZikNbAzYKP0YL1yvSDKE9p2l0b/r4iPtPfHbwdrj/aH3eB4QX7oZC
rhjgjpY488nZ0THiODPKtW9UCLNqxdhjE7RKjjKIqZuIj8w6ruYy17eT2vzdt9Ks93wbYIXmb0N+
38+86ggOqO7Vzgdo9Sb6CKqJwGd569aVMe1rZLhrpQ02KMEhIiQnL0MUHMRz6SKDkM1BHfW2CJsa
3KEOuVNQcFzN7VfIGaQGq6YXq5wnT5rfzQL3cxifyX5VyyJyk6pirw7SUNotrqnFP+ewYOONyncZ
uAHZ7JOOvzYei5TbDGWo/og+QlZlJBR8SLw4aAldzdIbTMclGhUCrNzSLCeI7nZ+YZPfs/OGO3a9
y0mBe7THCVJWeo4g+RRM1UWMte4pRBVbutSkvEqtP22ItB4BdDpSx0mYQj2rHerWFRF21aN94glH
wK8Y8k5luQnsKNJSixCrgGL+jLNRL4SkGYkmit1ENaSQH0EynLbizRJxdmD/2AlRmvDnPh32h/lz
go0eihie/xgLvsy1TvtIFXh6HPqw0ij6W69CsLP6eldqwl/+KcrPZMYC+2cRPFErinUu6il1R5qS
+qNJw0ofEns2oIUxFlmcA6YY0BHMQYaPG91IzNXT1R/gwF4eP+selP0TNEppjiNA+T2fQGwehw1g
DgvDtZBHIeN63B7RMnfZZowlY1gjzvpoZUkQ6ULrr2jaZhzPkh2YKliwhLIZYABNfOIizbj7Czw9
p4fFy0Y3ESaj3dOTSixh1cE1LQxslgl4RHjg2qznsl/VJtT26By9rjUVStWMZ85sdQaUvCc022C1
ATJnQSiYK2aHkX/lz/KB0lf3oW1n/lJ2aRX7iCsiqLBbgSb9I1Ym/ZDtjLGlwnSGL2J2H1SveksY
WOsOEwPkzwqL1WX2yqnWJRUTMVTodiBL3A7sr5dIUwghuqsyN2xxXVWlfYFNcBoMsE1va2Yqdn2b
GxHY3GzgRUdidRYOpFGMSWjDKPKidjvWd4i+ryyMjJT222BmfQYc7AfETcQTQUtbrT2tyMwzzAD4
ADO3WM/lac7WjXbXpeUWOD76Irn1cOJcI0AeGU98Wq5T/v0ZJFWMVi3AxYQPr2e26SBDA2SNqnZs
T0T+sEUyAGd7Hc8t2xzYujSWT50xWv5yYgJJexUQ4wsricwOi/6iuRD6z1Kodl85ryH761LxZJu0
CtWdwjP74PmvXQESOGOnaauXA+ohfanuPJtDh5wwVu1ErWLmGvlfCYRrBc8MAD7Gty6CI2F/5pJ0
3yVexvw1NybeFFYyh/55jwTFPx29XHNWJbBgP1GJakp8L+UyBfd3/PuZUImbjYCmeJBXkpdSgrXC
KaZeSUNWs16+esXNCe9uvRKCy1JeSYtPFo2ycIbwnzFp+DxPi1NMP1avzcXIUZm0WUa6saSm6ugf
FWVRrLxKwUqAh77DEJ/ZUPW8SejhyAKP95vJmfoVSvYWPhQsUUiBSTqqfwDOEhZ6E0GgL4T6xs+j
BWZtrFa0jwAiJPEGi7qfpsQyqGjMpBKllXGF9IBxeg79/8iNEsREBYS4rvbD23D+HArzfeCMpz+r
6Xpw9cDdVAqe/qV2YhAGUmSzIUv2kOcgcKPW0SEjXZAGrfowLkMqv3HVUP4+8tahnf+UqnPFhZ+H
vrs6aG985nOgcnXTIuky1QLFjmKjZ+Tx82gLO8V1VYfUlUfZIAWQYRFQGD9CsGB1+/hdyDbQrTiN
/6YXVdSoZenFt09rFIXsbf0RA9c9NTFcDDydIQvIb98GlmD4xFEaEMB1XCCoKndW7iye5Gz9nuVv
MSrauEv+EZ265xvL9VKkE6f0LAF+Y8kf2Tv0f/Va8/2NnoYGnb/Yem/Brr1cOHKCagEJCxiH8Dw7
7KV9UTyNKjsBg6zwFZqfscIDcfxyIvLmgs5CiF9bEbm4/BgmHNC18uzjRW3XpK5SNiPVU8h5qd52
K+MsnDAKDkN22zfLUDdjeyXRjdf0vJrxQ8mYHZAx/gGSJExQokt6ain29prwxpwnhdrmBCsBYhzK
98TjSnwowUioGvfk4e2FsVX2LjsPLAo1Fz+3OZFWhPxtHJ2zTsYbtrichtbpbLRXifbD3umYQ30Q
POgHI3U75UvGd8yyAW0V+5mQ5fa+dlPUs0I+jRakP+7KMZiowdvWe2Z7T7dJy1j35YP4prOCLWpE
G4338CA/xLIrEx0SJ/wQPk2eu6apExJ5IK2HK301Zbe4S9fpYxDtxOQ6NBwJsmss93a95cBtRbrI
dKOl32BlMLPKDBOBqiYK0z+u/tZ+Rpj/J/XrQ59HxaX7xWiyqGcfI1Fkn7oXWhtIKKN/jZmaFmG6
QLzQFiOC5IF45c3hy94zS4Ih/54ASSW0P1yf2OK6ubeO5Dv0rOYnkKnkxJV8ls6DMOkQSZUmoxsD
iu47JlVZErpPKuYEWzMMXpOqcTq/B0szrwTL0LoGb0wBKeDU+zPS7q+ARhSpKF3o1vNvBipSbOv/
I6O4oCNk//OC3sL9gqWkLRqOf2Y46BFeSUObT2E1pRd1NLm2POMDu/CoFKOySj/RILbymo4bfJ3H
DNBZdwm5fqwHQrIim4t8gh94eF/G/BQwkly1vzcFe1wQ/XKy/uyAFE2XhCURqXuKx+DMMMWSnZuE
llBM71YBLC5BAoqlpnbozWITZwZrzddbbEHKrbUTGYleWqNNgQMoTy53fT9RNkmfa1EzsN/gCkE5
u+DOzX7wHCaI8ARg9rNeetRRdT2HLjzT4hu6qws6NMRtRQukM8q9dEQz87XH+hha8KF2YU6jqI6R
fszsbY7ibh2O/N9Oxc2XXNHE2zHw4hBg/LQZ0C5kVfEQC+pMPxwCPmlOLzNcEGbgTV3hPGyYJreu
mlT82L2XwOra8izME1w7l61jG5mEiBkyWV1+6fc2epVz9jhDkrUgoggD9XmonS9Nd6X3uoWPWowK
M0fWjYEb6qm1FO09vlk662xAYkaqBcqsvHLny2x6gMTrtxydhrriYKItxs3mmkNv6uV6u8/C/Hjh
L4J1KSffKp8hL++VwDRtrlFMuKcZ46FfGUt+jc0NACPnzBdQwXYWoEt7gMfpdMwsCxo7cbHCY278
O5DKy4VfNRxcoeljHYLIJiJcImp2qxmC6wFd74duivrwgOOwzp8EC3PRO6wKmhnIQ1tUTgn3YRgW
swQhKkgXzsvvthOOAOcOA2NyyVND8ZU4Nv3PqZp+SgcVhDXMqbFbOMyZjhC9hKkVckj2NDTladQ5
pwp5Zx1voOHgibDmbvu3KtGDLWC0uqXJaXnKwhYeeSQaiCzlE5D4t3+d3i7g62gu7XmTnsUgI1Sc
8yd/n9RrducZ2wgjuuA0dpYlUuRx2IMQGJrgd9aOJqlVRgvWVPgQd0oKSOUuqjBsLVlmriqg7ZNj
ploUVsmRB4sWlQhfCU0RmkztMfN6aVJFxkb53ri+SdkTabP/xF2Hf0+ylT/AkcEnxe5JOBa38zbG
xulDYq3NoKSEcWfPG5SsqYipEPi1xLiF2KdsV4mJiQM1o54cqZ7S0sbRg/PxGVl1LiSc69BtJ/2r
LBKYgbsHqzBTm+9/4H2pBQiRqyBQ5sBuOweYc3k/VAEwKCxyeWXW1mF04RcOHTiwAqwt3hIRb4EZ
a8lKkw9OkWc3KidJW5MLZkAC5iaq2YTuIbNsuVN+D23wrrLQz2HI0od8dFxbFDGGQRUf+I3cgaIj
zgW8iVrYHsbQZLh4A6ziVV/JP8t834ySFe9EP38aB2F9AmNnh0TkE7LWwTEcrpmNtUcjJ4tt/CZN
J1XOnHCv2On6e6soRhDisZRl2gxMiDzWky82SriKI5VK0A8yQfuBki5MjFD5CaWlVI+O8lGoJ/XH
dsH7aUPLPFXBfwJPdjHj+Jl1+4z1QPgJR2I0cAxcSVEwtJOMqmvGXHQcgzwN+tfRN5vsZrRNpZYF
7WvcxihjKjPm1VzmS8RtfE9Hn92GGRecm8fuuHo6fO89pL635f9BvwkLYgha+WNMfKYaOkNFYR5A
i+EED2x/x5DC5wIjHON72Egk7NnNQ+dVIxOL+rJ4DBV9Cyq0NkuwSC95vkEKF9fgw81Dll7OA1tQ
8Bc7p8b6VVX6G0Qwy+K7SOpZUOpiExAoAE4X+4ik2Gzb5wOKO2aKXQqTUARz3eDI4k/U/XCvOtE+
3XUBCgfo78o56220VHaoxcP4dcOmStVEoMNyeVGqmWYbeDk0F9goq8TpzKn3WXaqFjOq+jAi37C+
2n/wQbu+WUJQRVV9ViXNUjRSaZd4+BEZioKF6ojvjLcTbPrr/QPy0CA2rgk/ayYG0RQnCPu8m+oC
Mdvu+AozDuuPDgJEHL0g3EntdUewL3vLIdCmnv/unmmGHmoJ8TPq1Nq6tU0HZTNl8mmJ9dP67eBb
9b7fb6akQg1+o/3MYgaKm134YUAqhq/swVEZDfo0cF/LKyUtJ2nrcvzzL26NzdwDLa4pb8uPMbM0
UfUsDPS/A8CdVbZUTZk1+qbuEOqdmoM+GuiJByWcNoE+JrvAsTDSj+chYrpxOf3m3jxa/+U6kuOQ
EAmSdIdhGKLzBoL5A7AC68O7x/ttFPHop3btCJh+5eXUG7gh31jzTqv4VuoFq2iB+v8WYEZYiqPg
RHM6uy/WV2wzdd+TFOVk4pYRqLSSHmnQWXUTZcFDUltC4Hw+bgiIHoha1Nxm9hHVS4cfqVsFShES
urniUwiyXm/PL4rqlZkW1NqlgSicStjoGsuROZpqvqBkf9IotNzyJY6a8qhj5cAhtO+TcmG5BBFF
mfehDIe7HZVJlhtmp2CKu4NHMEtuG+D2f7HGk0CzdkpHKHH0xJFI2XvUMRZo3xRaWXLjNScDeHFl
ouszk938qUnhvGHamgKUlCDipbRuMZsC3oZK1YXHFLOTYGGob78k6ISXNSiN63qW80U5gh+sUsva
LOtGJtBHxBbI9xHq42vPntjkSFoxWaKJaY3o3zYU+NK5qZLmTx8m+gW88hAqTwOXLt9t4tbf4L7h
aLhw1PZORCCNkDgL/gtnUlvSV08Z+Umq2Sk73ERXqxyBK58QydBsJfnaTXZrPCi5YIZg3ROncK8Z
smN6WW1Tf7M2u2SLt/wxV4CDL+zvCTKujaas7PXO9cD3eFOrCbPuuBqcC3xvxjBWNCzbBoI+FywD
cAiPECnwYrqkeLJEB9FJ/Tfu7osZ2NuiwbSOQDfsaxxM/diRw7nvcb5swloqlmvIVx8nl2LVgCXu
qt2c6RmDnUgp91xWY8l7CwSuMBXGFTDdB3PO28agXnBg9uXqwJn+TkFOToD4t2tTDPeBYDOtkW94
lnJIY9xkXd9Ik68X3TrjVG++II3FL/g1ebteK0FrhkLSi/DmAjGw8sIAyHONEgmU9ewHkUY94gzf
KU57nrZPT3R7vVhOnZXQEs5p8Opfj39drx81tjkdyEpqY+97meO/tInmZ+VyXYcJ3jrhYYUHDdln
jEYE/TjDipNDJjkwtKTlWADxzvbroJSRgJ5hIFbrD5Hh6zjF4s4Losda3iYXG6Z66VlKb64H/pdl
Tyd0jWBmLFSEFO6cNa2rnyjxQwQy2agOUseaZC0/2e4pt2wz2tSwJ8P5cii4625wCH4BUe9KADWq
sijBPX6jHxqAi6x9GT4bVMRXvZk5x59UG9OKa7xEzIvrW7Fizp4yE8NA8EBl2FGB+gpF+/vfYl++
KwWaCWwn/HdeYXZcy0WpPqwpRretaMpvEEsIq4Y72q6uOuY3Jn6jQlDuFyyROaQmCtLr9lteXDSC
IhJ0s4niq22pZSqpVC7s9S/G7/2XUm6n/yjpBbo0dBUO5YTjHOHoM0CiCVRUM11KwQlCPEhwULtI
vkezbCjZLUw2ivelGRew48lt4N9UPiBKYxQTmyg+Ec4LyW84r1SLCQB3RmBV+wxBvDOgYuvXKi2H
CgaA/hYEReS/JGZ4RjJl7x1Sq5eyJukzYe3ccZEKxEs+GmMLBS5sLdAIGlsEVXokWN100qmCts11
Z4boWtInnpl3tX4Q1jICuZ/bboMfteV4IAse+FV+0aMmO/TRoZL2PvV/X93dbdA8hhfn0cgG2zUw
6pSt3Z6eoBdWHzzgvfQTMXXOvWg3kviB3V+q82TuApp3efg4KIaOsONwvRfj77snTruFApsCrHRN
B14PVXgj5vE3LrP/5z2gVI35993F9ZaJkebkiLU9jCNLkzcnlpdfgPi3DnNO1yble/p3GJLbu85E
n/OgSSe+bn15Gn91L2ZBA0GkV/l/Pmt97xEszrSPdcXjSEGtbo8YzwDMPBRq7zRiJCGvZxy2dtXB
qkeWpfdMkodZAqyR238MDsfjP9I15kp0mabEIQdIbTTfr/rXBZCDR9sgD4szpFfLEvHQVOr7EZQ9
sZo9VgDb9X1EVN+MDS1E8BnFcop7kUrtXj4kLXW+USYAi8xhKxLOMi1R/2ok1hVAV6Ux3ThN/ZZo
3+GDVwcoPawosS4xq67ZWIgof36cGy1wLLBZ+6q1ywGw5jAho7hliPEVRreNhRHyXgzh1KhAOhAq
kJg3RiDg19g1Cs5+Vi7Q+Nh0xSlfy6WmXxuh+KfeeTRZabjnx0Rrzs8gz51ps92tRUR+4eV749dy
1SxfdKubIG6weJNjU/OecY5tsd/N5P70/B6+IuSYfPBfe5ev0hprcJ/AU+lfniGoyPxH0X1mN2H9
WwVqIRQ/Fss3Eivw7h++9GsVnZXHcvvqXTuZGakSoDDe8TX27o8OBBN0eBqr+nNnJCq12WMZczVQ
Yb0B410w7OdsoS2KdK0pXXpmUyeJ7W3BZK6JuHqSGPhMT7u+aWbe4JmJ+pTjMptZM0zLZSFl8TXY
QVuX17265yp6QYWAwXxlividZQ/P0ZYDJ9Wzub0fYz3NcsS6t9QRf2U4pTt5QyDIv6VBDO1OJUTA
McnnIb5fA0N8q93x+cAyHbZj91K4b39oiuuP7G6jP6X3lt0G5ekMKFNHgpnaLGgRvrXp4iJS0Lxw
osmRvKuNlXNxJLSaOYjsGnCjUhA3ylqkaLthQFGAQfmkF1EH6nSDs2Av3vFtj4pR+LeuFVePuTsf
vYpIqYiYJwSPXLlmBdV7ft0hTqA0XuzVJVU6ovHgvarbO8QBLZAMNWSMIJMkC0EAReuqC7vjJfIl
/cxg6nCZcU5dKGPD/OUeFov8iSQlFA/lNNj2iUz/PIlEMeO61Glu/Alt9Z9BNlt4gtdMV2pmUlv3
+P7MfZDkWcFq2QJHOb48MKIA9XxyoPY3qJiElEg3oWfYwKoqa7r29Hq1fgRQd7a1sWsWjhwc3IXR
2jIwkpCnl8JlQZ3Pp5JdNIyBmXJMMrXJQ8PQ+mWwT/aJbarOk+Hpv3J/XqxT883MORc6Hlz4kFV1
NvC4CB33PoKgB9d19klshHrupsLUBuyV4Jf/YcIRHIWieRFZEYH6MaFYxVNWFog0yTW0qNDftwtE
7tKpGC5R8Wwmtt3GtdI8vrK+8ioc7BRt+lFX81gQ2vn5m8lcYg9p/3u0DaFWlVkQFElhgw5n4wrL
EYZWSUSXMH+wRpXUqabKgkvrsY2gLfRNDC53g5C036ROw5QC/kTsxHwmRYMpp/tg3LnfcAzFhUPb
5bQs94qNNc0PFwFl/DV4vqVelazVB/ceq4tbRcR1i7GBf/ygbKTzfcn2jzg16i2cVG8xvyZudD5Y
nFUJcBBLWhhjt7aAvH4ViaezPvMqo591T1OaOB1X2Z/lCYsr7io9GTjooaCMziw02btLBc8uI+Vd
PCTQIcQlGVMWVL8cBZxQQQPamgqHKz4DUZlSH8l7XDkeXySJVK41zZyt8L5FM6O5BCDXTcjCLg8D
dMF/llXXd++Slgn51tuQFzotN3SVMnPvhswk0nSuk795laVd/ftiZPXBS4tdFJDlBFighXNi/i4l
lNjXzlJcKxi87k/l//9/UzE5YJcSinFBgQoYF8+GJyummWGUIxpmZ8eVx1+3XVZNMeSKn85B5pDn
hfSZt2dvgS+1l1gkkEILRcP1Ge8YyduUdGE1pWwvnvKhaUBYb+rDyT5mcgHd9S6g9YvQ5L7tcArF
DPOkbdNFHEgokRSbJFvuNG65i92pQo1WQjtQ/ooJ6NcuRML4xzLWwqWdVcDcOveUZblhtF78AjwI
lCpBkD835FUBcs/2M38N861U77Sn+ldmy5+K3q9hqrFXv50giF2d4Vw4qdvQfUYGu+3EaPCQPej9
56TVD95aivzyDiOj6KRIzp3svr+dHcPMC3bDrjzx4QUl4IjgTDMCpkzuQibn+2Xrj7IB3KgjXiNT
AgBNffCNLJAAE9WCYAuScQyyG9YPmPTtI0W41R1k9t4UHTWRobjayZZ6S2fiv9zFNz3GrKaAH4d6
pNu/u4xy8wpBGiT2LkjnP/HQnmS+c1UFREKHkCQ563P9vnpylBwGADQTAdV1v6eyswpgznScfyMk
KKhcUA10wVaHFsy/f5TX7bPWD6w9KI106BIY/AVc1ByOz7L1Tin6HF/pBPa8pzXmaf+5aEgAVe2J
QHGtWdilZseAab4zVQJPUAG1DKNaGEtEIsnkuXJhoGl9KGSJC78lBcyae/ZQJfdskXssRJZgpHUO
VZSAJQlYqHllKfAfnoy4vDARYGHZe1Qf5lXAP56IMX7yWo+HcC8KnKgU4vP6MFuvxNijLLLQTEMk
GoQmWimbpV3nhko6qoeQp8+4lqRipDMy77QjhWgK2zgQl0qOfnhJhG1GoOvDjcC8HgwcR1pM+t8N
YYRum9xyeGAHPlmttRyIb18+YzMXsUlf6Nw20BWcTFBA4CcQaAD3W3KLGDwgiTQARHF6KQL+8cOs
/hzvhS9zYn02bb/jXQp/VYMvJR+WjPfjYlzmuNg4dbrP+KxxNE8JB6Sv3sVW9PrCIfe2lI6KqYlz
O42mQc20l/zJRmrXxWBMPw/6bo+GbI6W84HS9Hrq3Pkjupj/qbz64cnmqCIg5xzG4hGyjXvKqlWp
anslf/mhzVNZgW7PbW7g0uGVJQPAg+8hZzqWnA5ZQ4p6HdL+y2nDvtvuiyzKEAtLwncecokct+Ck
tiYtTsBB4nrFkneDXBAdltC9fBLNpmV4XY/TEqfqpKDOcTLoRHq5QK0ikDcGFURUfCiP51FC2Pci
qEnXovNrBacqznKiaPN3gCh/XQt1mW7ItkKiqGvg+NX7k5WxObgsX/Edk4kryEjk+vWt53EiNimT
oi504oIDwl43CqkHGq3HmOMmvRwEudd9hoWoJSb2x7HawqPtMn5X1bmIw6IjXsijIkhyIK08nf6l
4G/PR5VMh0xNIKnsfFfYlCLI3hNWamCyTLZ1fJuE2yiFefGWkV8S3lYn2aZJ5cCLvHGXdDW+pU1B
8D/bacHqt4gtCYJSqZA/0LuMRjsjR2iL8T39ULRAmz4RpcRPQnziVjhjs1F0wsENl85m34kugoRB
sHKG5z1eQIDA2qPYPysrQQtQcRsxdqEiWB5OJyfGLnuhqPaDrTguPTKNzj9iUWtQUKKu1bJc5/T7
WHc+1q7UyKkGd0ajnl1bigIQKaJhXwVJA+7htAgE7CaRdU3e7sBlXGxA6Y93L2MQasM3OdIMSvOr
7Gc7dmaD3fGicNcP90aMDZOybTjbTP2SB/377kwKwNQnziaH2J1mS+ISdwVokBEYaH/l0M5tXpny
bl/ubgR1D7yMOhli9BOFExaG6v6ckcj6UVn/VZ4hglA/bA5khGwQCVdnYPNohJdYS2HKtO0LtyBS
3oIMLcl5iFHpWaXRNIAyD+onPvgSo/XJWmH4IOxmXIivCw35FKqcE8COJrX2bxd1YPOcSXRLCE6z
jQEDCddpaQRCgQbCOZdIGBAF1LFHPz3vSctSXQM1K1+9OE8ydRp1IZF+OP1/Or/aLoZ3Xnsj5FZj
DW25+4bGVVRONP+i2jcKNXz1LOFuz0JUwDlPcza2EQIn1lOpE7MoT/FgalFY3xKy0lUInFlGZkEO
+n4dDN4NQ8gG8b3asuPJQTNWqupPKSs4ZRjHaHe9bsnfvsKUd7ahgb3IZ7oJPXTQLquacDDIrEdm
gFkDDmb2vIkGsKTOJW3wqs31ah0JWSzKfosaQkfqlJMQT+SLbGiuW2YcQW34nLq0jGjggdCaU/dW
vY7LSp4u8a3tY1pklDEOrCbDthfgk/3zD2mUtb5J7XAwfkLF1p/hwZk5pP6zM2g4bvWFdddz8GpA
GFMK3EjDNi5sMlk/ZPg/yD+6RsBzppfGgsUmyKaNSPLTnjFBBMTgwb8nb3TclsLoitemM5Rz/Yd4
ahu7yP1usuoB7w6PcrheEyY5lv0jd9r6hRqRNqVrcZEgMKofKtehsr3FceCY1Bu8AyBo6zmpD4DA
xAf8NpmX5n6eil144D/gzlyzsCohx8ZrrwsU+00TGFwXzRKYRnpZNZc9Wjz5cmxPgjQyz+wtUZBV
/yqheldVgTNSkDiJx7ws7ERJYE87zWRySVyfWBex9hcLRpfDdaYI9dQkO/8IlSd2waK23I/lVA/M
qUZR7gpX9gCVcbtVRTCth67+XHBEgm8nPzzsLIdCwfrpJ2cHH6IDn96cqGd/vPZJxSBoPEo3Mnu4
X8W1CNAGpli35XELaoDbNRJ1R43fbM/byfofaAmOvTxmEKmGoOMDLLA7iCsO/2Yn2n5C7GnUEBJ+
JWmISAjTslmGzwfeMeIYBwPUKLJPcdT6lfKKT9kInFLebKFf9yGbMb8oeMBRIAmlwQDzjgDMIJw1
4Bxk+FfIe99sSQdU0/KU/rxUmts7xb/Ue1IsBs4j2tT/zKTgcaHPUA+uXSJMB1SGjU4GM/CVvuiH
HaxE/hFnvAHXLmtnMhOkhxutRQPQNvcu74XBoCAX0WpcGg/pQbiDvMV9LDBndd8pAuCz6EaevqhX
oA8ACgTfT4teOdWrd8sCtukRm5AK8xjbuF35cBAumP8rDmFrEggZ+n64ynAyRBxsgKWyD2noTBY2
vw9piCKQ2mUk+627lTKnzlSUkkmmlQR+MTR3HuZs6xGgBHOPPuiOeWpxnqvV12wbZm+kZuqqAdqe
zXq1X56dr0dT8/9MTm+9mHTlVxYfwiRekVFc594RUU5pjhmE404oyQ8ezDzIdDVu+jO5tIfhvUFV
FnGQCA4u/8wz0ZkJjO7JkCKNaWg1Z8/5VK9DCmhfcQYYFKWFd+M/LJy3EaDXsuNxBz9cppcLPbOc
PnNGQsfkwUo0f/O0Z3cElBtSN2i1ohk/bVAxVuBLS+NTvJfZ9yqEIXu8zltAauLVz12CW044wYy/
GWpToYgHd17EiOFAUEntLMo6uYYIEzoKz3ySbMCRNAGyUlD8HK/EERrfQ6xXRypZeHYKjoO0IA+n
OWD7rpS4b8xy+T5vniF0j7lCdBQ+Zz9kL2fIrDKn9VHSxs+xDSKqTKZpa6McWwh59MB6DtX9jvAc
XFAwO0xNrY5eGN96YEbTQj5C4oqQGJBcyEWe/N+jAd5L+R3ZlZkIca2V3kviPLetr6MNoh+w93f+
Hbck22/xqlCyJAguqpqP1feYFGQZHL+IfLRyNzs0zocN++MoGTP8Achum6SGmsprtwKZdKLYdQH8
i7R/5jGfC6IG4gLMqYOtjJ8e8xrL3OZkNXn2QDBzaDpiC5wNdLCPEAjVPBq2cBeqQ4i4YKsHOWGb
zgLqx+KTXcmcBtFD1qzTs3j8B1TSfVu12DqYhMF6OdleD7a19KeF0rgrPnoVE9U+IOUtpSgrwU9s
o+8ZtqRK9WpFVVLtPjcXL6WdsLh+eMEoroMR9V81oD0+Qmx0uhqfXl8IBFleSzN7fEclvIsdWU/s
7mmnVwQ2LyOkPBBE0uSIXAt9f6pQwIBcLtsmCtuWRUP3iGsnvl8kS2WaKMKVKUmSaMqHdck4mV9s
xzY6U/bcUz/SYOJZtxZatWef4zP/LpT7mk4dVjaK+NVJZ26FV0QtKvEbK3dc+7jI/uyjwjqTmiki
wCxJx8CAMWa5q9+XbOw/hZOd269uY4yvuAWquOcc0vBrO4e+LGvM/LHXc1kWZc8rHgImikjkh4y1
XEpmwXjGNoxvjzTMeGAVVmabDMz0wOIi1OSUiS2mpZvk2Tbngp1pqYkp9uPPHuXaZjEPXKiEyrGn
A3IypQlV13iRTnJxjjQ1ICZh7YwoXSMxEVd3L78BI4790fJ1OgO9ZfSQZF88L4khGGiG06rNFTY+
xBIcQnVSt+3y7mAQQ40+W2tfuGhwF0t73pBF0p7SWhwmhTKnJ1cTZBkXELKB5mjX/3Ealr+VaNsT
b5dPdgvgPr5N+g1jeczc8XgmRo4d17FUg6ykyitNsXE4dAjUAoiirFALc+tt3L9pCO/H8RX840cZ
zAv7WD/OaPGF5AYeXplmTSeyVSEf3/d8jCXbs7IvPrZ+DjcWu/PgMZwWgjyEqguZxj+g//Oo/8gH
4dDnBYN/9cca1bbrQnCUC6c7PMdBuE/m6KkiB+zXoQjpgKDA88RT7Xf6bs+IuYgneG8C6DC5SLw0
2vszhiNiNVDiVqyj1cIoqNqi58j5O9SCaC8OkCdNACzl7h5TVLVxXJ8JbANC44nD2wZMCKOTF4GA
bvU0ylD68N4MnVvyAwqbDclXcRwaB37aeMaXRzeV3DIABrzgfixiuRcpxJxg9kRjdEvx1C+qRm8e
i1z8ILVUxE7tFIsbPZXvXDZttXmqjjH7MWg7AwZavC+p5oajyXCNVCU5+8yvOadVQ1umBHaD7dMq
dVnJf7YcW6rJkIcAejWYCbkNwCyL7KSk63AeyKWLHj28wJQmebYImtWQ0ROMRNEklG+wbEkg2gK+
Ulv4YmczA1MKVNJDsOQnzGZdLTzRZBTU5zFTNwodyq48JSpiONBo7lMudIg4PIC69N+STSF70mCI
X3pd/LRK5oHkazNFRfo6FZm0ndUA8x0SglvkU0wH0/KpK67xO1i6K7nzX2Tt2bf49RdF2tn/sO1i
8lMo8BRG8Z1Uasa74l2wTRdeBO6Fd1qC9nXz9mDKh7X9QLCtVS/3qANDcats5tOmQJ3A78z83b4y
vBqhkw9904PGYMmcjmyNTdbWGW+uU8Etz0HC4Ko2jlDOCX2sIvDfGb/gDjipSLsBAnhlYSikkSRB
/vjv/uhLYFBLT+FWt6EN984MJafjM2NtdQw6w6HKdE5ce2O4JsmUU8GSmsYgi6hRdHCMEcvGLNEC
Ezj/5A1UtNiaDZ052ufjOdJjuZfWcdSdh0cAy2bQkIK2YSpRh2IDzLfpI+NDRYSYlzBjIHOxbJ7U
+9y+x1ZC9e6KPm7YkCWt8o+jXGQLdkgej3a3s1iDpKzE+LWL8Hy3LOob+1AZFewIAAsaIaV3O1B7
ewSqhgNdep6XugDDN2Th7B2ZXC0E7mNfLSeUiK7+Smn+PMii4byk1Q4VCos+hDk8ew11Dk9lIt0q
WScg3ljw4O2iRDWOZ+awPK/KUluA2q1yP19yh0KWANQ+sBCXuLZ5m1WHNmur5ltv6XK/DOTTNDof
Z4Xp2cuqeSYZHalc6dXgr9KG2k4gONy7gtFq5D1D62VD87iK2IL4q3lWsfVUc3Bf7Xyxwu4IUi7T
NJ84zh1GpMVTL+Dm02TUAtEZeXJkXK/Vi+PXoGP7xjuGNHmXsK+PWtaHq1BHwk0C+GqF9PxUlYNM
NSFGr3vjGBRUNZDxkgtvJq3s935XuqIMGJ85fhhmilKXA2ULuk9vWg9ir+eL8IEXu7MoTUew9G8z
TM9RaioRti01KrsA59gMk/xQooTWZWxDxEIFqxi5qzZY8Xo8icRWxyKrYaFbp4vhgU683bFAsVOP
z7jiExe1gQ2vwp9itNWTk0xfr7MzwHRKkrmKSUpFa7BbfgYPI339znRBOOkc1cxTj2Td0bfDSqqh
extI+Bno2zRUa8iYz8bBzJpFZxit8VEOmVCUNnPWwym+1oInTosFObDsMHKbMPdqeLz0KDxg3Z1/
IjrRXgAMIUeD1lMn73vREpv67f4A7uBOV0wEmt0DsRBykGKqcB9MNsdma7w5g2pKl2/hCs63Zwig
iWZOQrHMNdIey/ZjmOs0YdWmsmt/AvnafA1ppiuiuv53CP63dviCzb1EhcMHk8xBBl3OCwxdjjOk
nz1Qm2s0KNGi9mo+bp8OPloF5NDDTQG9quUVc+0Z3R2KisItTacND5kk7CqTk7dH6ZbtFWywbhcD
jSYlIZLpGQuvUpYB71pfTj/280mQ8diJXOSdeVlx4oLztQ+ES4T1KbnGJYGSlHlMUcmVvBhrLW5m
7du3mWBIHdW7EPgqldju65pRzO9d+f5Qo3/NwDuKcDWKRZFnDlxEF6zBJ4BnDdz2Kly4BVlvG7pG
dS/tFW1VaFeVhIJNDVnwrWmNPRuYHJ1jvkdKu3hNG3ir/qkoNbJfKrWGnz6ZPuWMBf+Ue33L9MSq
15856/H/+MLjaf4rKyHG3RiyyjcrXRimWxtSSdBLHN5VzzbCC3lBiX1Jva1ThqPdcwt+1eYjYYFX
FGygXM2J2HDlxwmgQCvLAocAOnsuhHCUX68Ybk9yBTTyeyZZyyqMhnggM//MSgS0elXjRahuvT1o
5OBU8nXKZfymhpe70L7I4ZvdhVzPcfesFsoEyKEFRO4nA3d7KurY4v3WqgI7t76LrKcRalh7BHIv
9tD1I/WPFfQ7Eglj8x8bWH+oH7jiicf2edXmOOLdwFGrhm3R7iK8t+U44e9eBTr29pt2NjbsDmqr
BhD74I4jDP7PblYHW1xm+eRF47GCsDEplGBZHINzNpHE/wnPJemdpfdeLPbSVTBVMXTGtUKi8nem
Qsz3L05KJMDNVvAt2SY16obtT+zUwcMi0mjOKlTqEIIrjIzvNBE5frhoVm8oga75JSo4ZJND7yJu
UZMcwgyT6LUSzCy2mykDgCf6bQqDKSvlNtOGqFLjC/sKkAxxrHcffi3JYrI2lsKjIZnRN6hKmpXq
SH1qN1nl+QjyJkKp5FLkFmqKRhOyJqKa8N5kodGh1OGfQ+A/bT68JvS/crX70XUI8Y0Vb8r+Rb4u
9ESyOSuSJyWfFo6CxB6bkuya568yAluaYiE54AiWOi0GWJ6x2LZtM1PJ5LmUFD8RzAG8c+o54PDH
cy8FbVZEb0mlCqo/ET2RCBkCLG3dxAaO2OfmuyciWzkoknNNQ7jdOx7q1FLmNpCHuNIbWaDXx+/d
HHxKx5UDcvBc2ZfUhgUdSnW/SHESbDZ+rvCK3S3Zqliu3W/DZAhgNCZ2WhfmANdF1342HRUHiS0T
DKwi7vhN+ctXDGDVj/pL9o6X9Q+3vhI2MwledG5NCJJgZsmTXjT3vidQ7QPg7jStX64sbLQWe5p+
2a7kaz6yTgohx8tpKxWgNblwiITAzNNnTLb4zRVL1YAYqd10OE2Yr12QSfwmaJ/gI7nAeMPHebcT
oxboyynzATW9F0dztHTqGjfyRVNUCKevaEQyCDR6nMdhHgQifPHUxlUU62QoB8+7Fyi8/Fwdn1LX
g1uL7GpgwP9RnqKYSCM/cT8gmi5olIoq2S6LPaPvE59H/99IlqqpIcL/IYe78GbuUetNKwxnYazk
u6xxhjsBO6dyoUv3edq9yKfwmE27L0qHZ99dRJvhdlSbsT50pNXTY/m8kuaFPZNTrTn6Ktpf47cx
PXrI4r2Won6KySQZx7OBgBfbUlvDQBYH8nnWgBj37wvkmCb7N2qWHSPxnupnuVHmrwmvZWmUAuCD
6VCV4cG/qGoy3ZF2CMAuEsAQ6JNJ8CdBku9QWN8p7uy8o7DAFQLxhcQ2Y4yRxdd7gQyFHg0riEz3
+/4pN/PgEAoEckz+gYvZNqmDtCn/CQy1GBZSzjzYjR1tVsUMZPjBhqCyBq5P4ILxBUt3h4OkeJTX
VtcoM9P9WZROQRNH0Gg/CK61PTrkzb4A33CzCJjvOCOOMioyBhn/xeFqawgZusqaU/nRthwTtO2m
gevGGNyhPP6CVai3NFdDAAfVWZ1FgXp0b3bPu0lSDTf2LXAPLqhQjXpzP/cx9Bn1OxPAvQXerZDD
9HEC12iWOctXO1+OlghoBwfCJitrP6tS7TU0qiibWvYEEk/47JT3iWJZRy33tB/3aZ9l9h9I9zfD
ONIPWA2nlSURjqGx1cc/8kDn+Nz8zLHxECQrzpdfgF/TWOXtwjGZsgIbf0IE8o9Sqi0wCNDl3tta
Fnc8SqQVE6RUZbGbQe3Eifw7Ust8qBZJw03MEPaICNc6yQj38YPc/Bng+pqrZipfZujQE9Ytx/d4
wYUvmpjTmph5fb82usi2egsRkBEabNq9WSj7dKpSkZ8J4FmV7k5zWVIo0aLwjalpmTXN98gqpS+i
8xdJ4q/q4Yz8tS8qjeec5KDQksxSpdXMtcjL/n+BOuVhlgPGCGmfEPCG6msmvL2jJkL3p7nYjQAS
D/EkYOXM1AL/+FkSoM0ESOlpHdhctaCbYhbFqHQFcYPsKkxUtIpP6vpZaIkgjK5fc0up0t4YliIJ
+sF3tH8uV/EqrwxyoGdoptXKzihoeLg7Udj9UDLD235GpEfZy8INnSqYl8tf6ierGk6vQDbmktQZ
/2O1CPfjB0/ECfeRZPnPqh9ousrhBa6NjQ0h5fFY+3FyvcIYglU6hR98X0fDfUqmsG7vQq3Th8i2
AesNfTOESz9T/N/lYg0qeAradePmLmISMBgxDwM4nJVzqQjEdsyi41iTkoVszH//19fTtGNYd/Oo
qUOGA/wY5EmfZhYNoO7lNsIdmEYZkKcoH0o/mokUnNsXAEvIq5E1e3EWr1q3CmZ7LkJNVAjLp5ER
a3Lwqys4ghoUh9/FWjVuMSLY8vlFpZCCgMNCFYzcTn3IV+7oHHe/YwZbvjKQHm/oQAT1UPBhAeMV
Bo2YBDlNLD4Q4UBvSlH265YZG9UGiW5zpccgR/LxoNjN6fkUhclE/ANxSRrzPB+vi123ZSP0YG3Q
2Kqe7hg/KOu682ucGt+Z9U4i1FFXrzUG0V2727D2OC6wmyuoFYOtLEnhJh9mtR6KXFOiqPgIMedY
ZLGZMQmcELa9kmjDHop9Yo1LpxeyaN6HZjDJRdQfjjROPoBbVAzFvL6RRlqrLfzd4GXfPx4bXuTM
UqtdTD4wKrcDL3/rv3X8iyTzl8uBNezDbFdQf6gxu5yY/QbS+QDnJ3mrWDe83mQGrnXe4HJO0YAP
p0Eo75xBCaljK2KejD6yBov2LGk16uF85VGb26TVbHS120bYR8E9RSZlEtFdcxLE8jW0aBM5LUXp
ds1vpKLzLvk9a7eu9mWKCKBIqyj4SJCCng8HRA2e1IKsjfRYawCLYPyuhrlXj/8bZTeSGwEPipT8
ikp0pZ8HD6qIF5nnr4zqf2Dl2Jc6NJ9v4kbad5AZVlfKamPBcjrFi2w0MbYFORemIdJN++f9P/hH
ctAyjM8oUoleR3S2ZkXiFYVVaA31m6U3/z+EdDsmJPqKRWqgnMUKarNkty6L7jqBOUc38RmiBuzW
wV/BaRQ3u+dAxW2HQ0Vm6DOEt/WPf5NooyqH9DkQwlGnZk6GlDt1rhWl00fBqAEtaJ/egWfBmbKl
0kRtR6WgCsd9ZbUVLkr8nqLL/tT8RkADzWbukGlbW5kKyhkJCuOpFtwQRym5UDRIgytxOO3Bnwqg
QyllBcy0Cl93eJvvWZ05N3c/lHEJKsUgDQ7TyYSSZD2arlEWZH/1D6AQ1GsCS/crn/N3zhPwKDJH
P65qNpZ8XSazdfeE1zYHvboVGwdGVVcUbi0MjltiB174+sOWkYriR8x7j7NWAHKx+L5V0kHUHdqW
Rd/MkJodg8XKFZP0wYWhNSalC1/2C5rXhGo+5MM9/WYoSPcsL6OfrTCjNNxFYweo9x99VL7KpqUk
EnV76oCp9YpsQKpqvxTDMB0qSDwj7tKNLlHfdH20+RXSE3rqPQRRx0ZYLvo6Yomxk6gt0OWqzkzl
1o2XhG0ITAaBEPwYh5dz+XHJgeNFBzvUhqXKvMr5epuOu3WQYvy4h8Sg0iAmzG64yBmMwuSIQMSM
5bxIZEPdsOg1nb63Y6VwYGWQ/0yiqQ6ivO/B9RAjRDCLjy3kknxs3n69nwhgIl5NsWFFeP5nOIbJ
IAPndFYqVYdWSZfX7XIs7BkIJpga7QboW2wgTGN6J63IYIf5XvQtWAWJpV4qnpPtQu8xIc41Iwp0
r/f7b8Nr2eoxZUl3lr8ypNq6HvkWXmrL92Kq2o+6yfVnRbuQB0Mn9uf1295xgZFm1xfbvEMCPlWe
mDsSbKRcYOa0GxBHhJqId6XHoyPhYQYaMexG05YoDoF9RICJZvjU3T815tR/hM/rcitL211A630c
0MXmfLW2+EW4XV7vzDM16LiJP2Z13oocUBTx0FLniARb2XrxQk+g2A1ccn67gWGfCKMcKex0nnsK
+vF12jB987I7hl1IMCMPd8wNEntUugJ0jBprlLU2/5KlZ1tjJIPhMXhrMUym385E/hlaHcU0E1L0
A4/7Pmyq48Imk3UHvlIgRvAZfQyQylQsONSrjDFNFfHaz3NsWUI+JAPZIh8t933PKTzPlrBju4ke
m7olnd8YOSQB3dq4NXl0M4fsO1kwlqTo2VV1Idp1vzVz5UEmTef9rjuMVYpXyBMuU5NYWPyGuJ9U
LaMJXNrqlK4wS52G1IAeltTP4FFjBaDnHmh5s656GoS+3K4TRXxWW6p0gBAcsMswDKZohi+y7wfS
lc8MoUkIPz2PpBlUyofxUpkeZtodSe2DHmm4wBKeOd8GZyOnb5QpQNxOqwseDVbq65+Syxm1SW9h
KQt5nKyn+iGt/piregJKUAMX21bGuf7/vQIE9KWbOLxEihcz1jociFnZv6VtxeTpCjDVipTBNr+7
How2QzS08ibff6ph9IeQca8iGCnY4IDsUBUFAudytKLYCK02gZVJ0IO1qoUHDMObvJDsKgDJryjU
YAY9GZU+7MmKijdT1qT9gLcg/wKQT/Po1YLwLpTA950eKg3DwVdP7D3GIUlIrFZKJVDOpEnvb3WX
9PjceMclmNm9HUIcbyplw6zQ0oWLPBdSktKJZJI761pxVaHbMzNLjbFWhLwuIrD8uxv1BnBZevHK
E6C94cYG1xOOadTQW1ji5uwl45g4i+qKcOT2IjrYRArz7CV7PDVtIJ0soeGqyc2UhOl0k7d6Ae4/
LV7xLVSDUIXeu7aIlHtB5YAkSVAaMy6nbPHgU7CZYyKQ+1KMNmmR0puVVKSSiYkHRLcbEOg4Dp2C
pLYyAr2G3X+TAi6vCvOjv2AEr+fLiEZApP35fDihLML+ejm+n4UfTA6lYkPYF492QSk2n5GltDNR
WPParAzytACoSLzxnul4o3q7EbOGpShT2KDtVqWEFAui3gI5t+z6ELNCRAHu72TMAuPJiUCNbsM9
Zb8+iABwK7AwZ15OdE1nBR8DjaW4xKQNMPS8SDMbdi9638kXDhTT14P3vWzSd6xEu5R2zilIBdGy
ORyEGryKPey33MObwkSF0EwR1/38aDCxO7dLovkubzkn2ZRL1HBnkGpSv9HcUNURRKbbMiQxySO5
fcgNfuuj/lcC7OeNgR7yCSxX6VWSIb9r/8UsLEY/Ial6a8vfewWLNMhO/zL8mba6vuTFMRKQnRFd
cisdkMUvmxlJi3Q81YFgT/8Fa/6jNqW/bIA4CaiX+h54WAcxGO1UlRT7VVZitdwww6vQP5mW4avB
b0WfPaRzrksSnhGJltNJs5OTQjj8fbhgazhSnNqUTnMCTjdAujJT+FwDUQSX1zKYguB35CBLmlBB
P1YSMu74jEHyS6H/Vy7VcS/RfiwCkkMjKuXIzCpq4uxwkQszne2sCJ6MpsIU5cOXQvH5l1KFWVrS
x5itYlJohtN5s/YI9Jji/Wkf8K0LS7SfU4a1Is08WbFywxyL/cfos237VdIMu5UKMY+8dudywLEB
/xBaKqMiQtYSteb9BuM8ycuqGV+ObCih5ORc1yQ/GZLI8aI2qkQwIkiJ6jTtvRAgSmLGDXybrul0
paJUHNsE3dej0crgL0n4F5nJRuGyuOa161nyxbr9seZ+eVduPDJJBNd4Iw9SSdm8B5H9jYDuTRXS
wKn6XqkGbjJKsv1TDwzIqxW1aNcTU1k4+b1DNFqrDSFdh/A1W3hrDZwWZ65P8Cay3ZF4F8Uw9DM3
6O4YXbGS6aOxU9fWHvfXGywS4S9zZdP0jAHuAL2Tg6XaaDBW9N0jokduSEnf9bh1nLykh3IjYgRJ
5x2F8m1pm/hEljAjLbuyppg1u74aktLnIOkO+dnR9PeHgfsTK5H91w3F+chTh625AMaVVhCOgoEp
vArqazfLj8YvaB94pWZz/HIc0kCr2Qb+E6dzFbsg7G77E9o9svDnIeeXcrVJPzef1rXFSiTeVpNE
3hKXT1ysrhzs9eZTiM3HGR+1J5BHYE8rniDvIRWI8fOMR2BQc1l5UN+ZmBQrpK2KCBtOYjf95N/p
76uDNBCpYJoJjr9+0rp8GwAcfieAvbzcjTxqYL70yy13s2wNXkh0UHdnLIR/4i7h+i7FUmUUWhO2
Q6qmDu3076etuujjT8PG/t6/G118hMdBlx1Jk9i5rsubFJFforXHfAmeGK4k5NdCJxH+Wj1gnit7
ivGObLgGa7BWH4tJ/0kJJ3oYZ7t1KWD5N+jsh1McGDcT/nkEfOLEX48aC2hNCFgQnaqYk50QIslk
sWclwFOtW8CbYLMkuGUCAVYI4KEkK8zlb4aS+hvUvwrJQItnoJKS45Kbhu4HTCDOlE7dl29vtm3v
e+LNGBd2NQF/3+XcwqR7BK54iIBvF+brdQaHhiWqX2lq1nt4A6RT05YR+vcUSLzE8aHCw9ceXHj6
WvHZOv+oIMKvu7drwBi5wOTUAV3cR7K2IKFxFjr7mXDw2LqXPtqwf44G091+jP5HwWWNJNpWOJHt
l9FPVlZ2yorg6imkLHW+bkpzgcR7qcxM+VBZMv3mKdlplXayiRyjiTO7PyfLB5RGyD6jN/oThHOt
u7LWW0uLtzCCRrODwaaJ7MnLtHt5VrOB9RCIRqtJSa+X4yYMCBs+h6cbDwf2bEUIH+kQDtl4XR6W
SMQs5ZTSFBeSQ9S7bZQ3Qo4rLOKAW6tCU2YWIEK6bPXRzkc6J2FTrsJhsLVtxSbRHrfp9ifVqv8b
hupK6i3YLh+lvEMJ+P3aTvd0TOI/IwnLBYXv1ZV0UMPh9lMAzIyVN9bm0Uwa6gYI6aHV3Ha1VYbO
xot50ycdyB2pHzrzYJh6CEODl24bVVntHhgQn3HqRRFLoDiuqOdBtkxzpmTBS+pqVoWARN4xSfGK
yo6N89R11psw5dj+V1XnaqC7OGHuWt7y/Njj5+/m51SoOEPgaW+iG3Dae8riv14XEwLHMW3nyvYJ
w5chv/hhY5GTJwNw+3Z91gG91Y1+6aTEeOEE6Bo1FqGb29hUXu+85liDyqutV+qUQQb9/5bZXU/q
azCf0RGb4diACRcc/Sm91gDtPuNXV2WZ5xiiHvtCMD/Tu8aYAdKFjwR7NER4rmFmgGXHfWJk7j6E
pAsOLHXybPzNATFykMmoG/JfEMTtb6wyPbujYHFUMrM3QIKqr5e+Y2g00OgX9qbCKQqa3m9ikBai
VzVOhorNrBSbshHeWcyGcf0s8eA+HwvkaObyNZioD71MbvUQUFleyO2ZmzFoVNYiF6dJJRYxiztP
C3+jkaZMFOBcMiCPdU6G2kVJ6DjXV3smc4/ZsDNaAxjT2xz0yQaSLxPb9kAy/gc8NHfH67MvS7sG
S5TSTqUEoqH7ugqQ6l/nOg2Bm/OlczDYsTXSSvnEtszuvDFn2i4yKmHOs4grb87Tp4p2VkS1hc9q
6xqOZppoqHGutp1tDE+Ffo8CFXCw11Ixod0hYR8SEKCEnWlzHj/j0L4vuAzAszhQkmMHcqi0ThuB
vdR6jfx7pm+jnAh98mlZW4MONylv7OLJE7DYC0m0UH261wCroXHk+vzdXv61fh02knai+RAUWGxz
y2rfURbkSYJ8bRAKEWvhb6ze1x07eao/twt72di1I61p+C2TkDBBPbADXOaI9FXlK8AAqWCs6lbr
6W+1pU8/4rV3FM183tg+BT+NJosDPiSO/9CzgqXxBQvYPDJQssoUtb930MnsvIGHXL3illkldOWm
HWCLzUdZOHGE5MZCWdci/sxhfyaaN0taqdO24ObV/+2f1nAao3EIeto0dqGbQfoOeLX8AAeVZcc3
Obt6x3JHuyzbr3ZxLDbjV2R5sPqhVGpi4gI8hOZsshD1CfXew5xXleesx54KTkVb4IEVWndXGpv1
J8yY+9DBoTkDqPj8akXFKf5W4uOa4xyST7QSgQc7AIgqIiK1sYNSm6tSiGdjBZDIMO5loXeeRCW5
GiV9IJT/hQ+NeW/m2bM7xq7XR0j4sbITKkVvPgK1ZmIqV8hva8K6S2PlYOiIGrNjU2FMNwB9rh5Y
mzLSUStQLZbcwM2s6W9jdpDQo5S7AsV2fRrL44dqhSgT5xj2nDUmoTDjrGoIWBFv+ijwH5ya80AU
J0MGyAanW7UvzYtW99n2aIMjuJK89oyN7aS5ZdSDX+g8IzdxqjYjbTIIT0u4xNrvMCGTa292EbUU
HtsKZhz6X6UZEI75G7knAjnBVeqbuDOJjvAKVXNanB7dMEX8iOr5AK9fUM4Z4I+KUuI/qBpE5Oux
nJH590gUHllRomBWeT7tBkWQfcbjSwfcvzXNYGxLmaDCbSfkGU3nf+ubBSEU2y3DOM0GvlFCTPfP
NIRc0jhFAd18yZHKc7rZVlrBO3h+3VVO1Yvm+hQYmi/YWaR+/YpVHc4wS6Zz1m4tbmu85HzNJMnl
Xm0zcVl6zlugcrWlvihSvfX94y7h1vYCYQ3LcE/Xzr2pLYeUyZuojMGo7BscVWiQqVt6EJ5cQfwL
PmYL+26JJF8dRdfKIaBp6LTTNtIe8ZKNFBfnZmOyTXVdHelSxjPeV9XpTVKa9mt/9tGunrktBVpV
LTrwr130jlF5LhjGRaXH0aW7SZcvT7u2wmKZY7NcfM/T+npK/dqkDGpphSxljH8nofiKG+sa00xF
2w+8i4m97Ob1sPPrtKzXqySB2BbM9Vvj+/Sns+0ll+SguwJ7xymavxvYzrJkkPK54jP9jKwUe23e
HVhsX1tWetxWJT3Csz2eiZCeMT9LAkZhaKATIlgFGEmtQ/Fhvn6hf4yROGxEXSQjGBjU7OfDOmi1
ym3wjVDYDaP18x44/Db/XMANAQsboLdiF113U1xFRh+NiYCC+tpq/VJbreFGn1m6wjPxsBBTaO0j
PtH/Uad378HnqQzc/oKB8Rnfh1mtFRMFiv8BUANdOkQi34t5J2idmVLaf/R6BV3+8n6ElXFTbfNf
C4vLZP4oCMGG6pcNdcEetjAKA3Y1nECtHQdIwlXSmDTpuBFAnx3So+VKzvFEeRIY8h0Ki38Ke6dp
9kXnu/W3suOagq4V95Gu3OqLIWNNMSZ2GHeNyZfH6FDJ6Vi+a6B5YlyCvAjACEnsJRKoIQgvKiwH
qH0soa+gMsatlO6c9aX/EAnKyLSllj3aLvOnxjbeMNFOzjmDHFZK/UIWhCnAtkU40Y/fCeehJMsS
IorRTDHPy6+ahgxvNgfKz/9ArcTao9bTrWr1P94zMkQ02cNwHdIItZodkwB9AeQkKfqX6ORVMeqq
5L8zTVcUVhu3cOwiIRb5DtpdXnobTtF9NBXj9xlO+9EOZm0aNEdOBxLZkXEoryR0t1FCWzJ4x8XE
VRajqEjsgv3vXCyxFmFirjHZg38qdnynQIKxYASico3fYTTc9m+L7P42LqtVfAbqhuDEVph6qlrt
LnUHF1mmshjeWZHIF7LgrV+I88Kj8gjTNaaEI/6mvfu+Y3taaphPqPMPoJWRoJWsDfFX3wGBV9xH
0xsfUgYQpjLMUo+EeextrI7VaFqxRLpEPUXjTsxNkQUK4GposM7cUiICExRETKFuodUPad0+tP2n
XS1mC30io4AzQ3UeAiLYOAeB7X7bYDnCTLq+HyGfZxcPnkpxhqrye6dTC/rpwIvc/SvQfUGpPqMw
gXC1HPzZf8YCPLL2yB0TeAt+t4qmGF8X0ZvzKlHri6Y/QC0mzIL1WewIIsCw1DMTNIz6ghV62o9o
JJvc7lCUylW52FkUFlnDTCryA7j0Hzq7ijuAbkO75T46+N8JY9PEaihnwFCNx7lAEqj/7mIBFUIp
QP1XHz2EraoBMijIruz8ax2aEMkYmIqv32e/rh/BBOUf6SXA5+wEmX5PGKTAryGZRhDbb/ljh+7k
telG5hg0vBQIiJGAHzBeadJMx6mUGmvIJjDXzh1ktCFXWdvhgK2mn2g+bIsakcHX8lxnLuvfF9OU
aSsc3w3REm7OkibsE69diX3dUofsuWeWUmQEGX6ltI3XIsNrG8OKf7ekZf6Z5Zz/vy97zOnYtzoo
OUDu3Pta+EmXhYuO3DQLgUqJUXoNXkipx7inB/9bH/NtPjuUbCMgbKC7q8N/K5Um614R1Wl9C3Tt
q3zinWxHVpmBjnqqHPJlkJkrPdoBJNaATEKWr+2ws/I1YDJ3UzlNditDDR/fJtA2om68pOEDcoPn
a/rbagAXFJXgOMQxT/DD5LQ+kP7bcDNQ8t6aG37NNQ0mnUS5Z8rgdEgS8rueXHT6BxrjeHmuqsWA
Y2PnEb9Qf/lh6/EJqN5KGwVrKw7EYSqinK2JusfTWCIg2Yr9CwvqnI0NyiAEFjAro69MulygnPLY
6JhmImujg/1kuCgWq+9FATmV+2lj6NeZxdNc0A/L9Y8XNlW8YEHXniDX3Q2/ctGI5w/JghUlUCCQ
aAsPoLwsO8MCqoV0JIRrbEh8dITwQ7nr+xXLvANJLmNWf920HJcxYYRKXkTDfq08py3hbIfJBo1G
2GJiXjpzxwcZX6UXZyfb6b17nX4DZH4jIdVq9Q4uJoppor0DC4WX0aUoNeDhn0Cil16zcefmFgeq
MPan69IZlk8Ic+Rj/32pRUzMeD+gf/Y9LwC6MDcI/3YREk0IC0zdkTXQ+JH2J7klDjqWvXaxRueV
59EZF31gjX0mw+3W/0WkeAZR4b0Z8HzbYS5+ebgixvF0D3Ns7YVg5XVCFsbUJH+S7iRpJfbwItA4
Dnx3UXuN7orveEz7eFUa5qN2gCwNdUQaosDJDcmL0lK1xMlf7R0aNsfC8+lyBB1VIok/cr2+KaLg
voIXw5OT3PZen8z4nr6QQFElaoQop5VXeRKGhgQx6sjlu6rQfJZtayUvyoWX62EKenJUZsa4FMgT
VtfY+egYpW0fc3UtUVBlBtypsEg0ke3Ch4t2qtkp6k9sSl55Kf8raW3wdULN4qY77TQN86XiGzTP
/AoCL75wkEMpGGPpJm8LQ1ayd7K/iaaVy7/QLq2rLYbzaCr0udAxa/g4RRp9a/zmM8Dy0/+7nDal
1zCtf6wQpZZXGez3vFOyhq7xpaoBwbF0MwPfNu+rXlnd4RByCWXZLrX0rr9kQcmmG/QdVIQGAcrL
rJinGg1NlVcOJfvLPMTN3GBBEoF2bT+4NvCry1802iBkpuHmfENflotkj0f3aS2zM7cvxcXdzZIq
qJQ2gN+s08WRUxn03DMhhuUsXXqjI/bGMpmaY2JKGcOcqpUZtrdxPvLVtJiJmdsOWdx6jaWDhxd5
mrbiwuCD029luV/xAEisqd8mpxKxL5gwQxRjAPfVT5Y1ejk7qIdj7x8cHkYepDFtEB9LW+SQeEt8
rpUfgbBmnWFvULe3NIIUd+nWAADT6ezDFnP8BQqr8MT2gBb4b0y4/evj8R+x87IQDMDL4CSeIgD4
bUUt+EyBZY8I25k1i1IWNACKcJfO9h94VuuEm+qkwZDP022UhbhGNON+euo/R2TReWEpzRLjx1qU
H84+mFwqFFB1ESknrTuQYzsS7vklGjw6hfIl8jml+TnoCvrVH6EeQkz3ie7Ukyuxfzs0GXUTYnSi
ge7lioVvIV2AsI42ksc5Nq1628wNPEmiRRcRkCBWmdfvdQEXQHfM5T1lRtDi0OF4IMxTS+Pec756
+a2DucQMaKPrhsEhs4vzSGrNBWMIPqAPotuFjMkNU2uA8uP9arBvb3UKkqM6tHIqnom6kVkcGOMN
cwQPWOxNeFw5rXrexwV8RK6P0qBy0zh3+JJDDcG5x0qsh2W9QeE1niGWFU//hKr05Iob1GnOGG9I
LQTg3a76Q12zfuUfLBrIx0SK3GaEqph3sZFEMVTDRB5x0zsrgcf5aJfEP/WXBGrYPV76ZSgqResd
GggByAGY+3tOxmg+ZrF+fRkf3dl78r5bJjzZ3YsIfwnTmMrw64atPej8zdbipSs03TmT3JS7YoIl
AjvUs/KMPA2nzUeMKws53QAiENl0TroMn0VDF5MyJvMqOyF8WjbxeVbA4sAQ1jbdVh8VLFL3QHlz
MXLgd+j5U4FPg75mpfLlqtfLZN/Zpn//KJ/IPs+YhJFFbjA44JSYYRXWv27zX/t1CVUA2MEb8cCw
9IFyhckVSOlux+Un0Og356KKXRpKGDYEg0/21yvAjM3l0O/F2U2ICgIF1jlNt3EtsUp/fQoLk+KH
rxIY6Vh5jIJnZKzDp/+FXTwYxS0S93sFu0vbJhlpynfdMfoOpnYqgJk+0G2yJJCmvB6kCk3TcAGt
ghidovAy2na5FWdr5IHTyAbJ/mnfOLflnFGO762+JZ+mbr8fFcDnPKvhSTYaQGzq0rK3H+Uua7st
I+MaF+G5UxSeJo38uQhzl0u6iGF2oz7erPgvmu+BBAnIcDqpc6Ae/L3cdI1G/enO7Xa9M5glmzs1
+WAZriDP2JT+r3jnNnw1hrsZI9FKWzRDdw+77FLsVSEarJ+rTQIupSuK0oLhZZ3UJWzlQ6AY0jXH
uOphqIlXAG4a9aDzo18a/AkW965GmoYjSltBpIx26MFaSvXYOq4FP2hFmWbXmTcro3a93WGaHe3h
ppra6PgOOjfzyy2KKvBdz3t9n38DFdBjeiNdXgfYRlVPh7kSOenNKLOuBhTL6q/SARKr+rwFfgGS
hGIlsSMEdfMIPwjL+Y0+etUsAJAdQuJWQlnw9BLbnkZ96fxArA4X1yj8OIpHgyVUSaT7lD42Tj0C
gmrEqSnNXEAPmDb+7L5w7b68USbplAReQuNp76DbOiaJ1mQ7Q/YndYjEVl18VZ0fc5gUJ5d7m3RZ
8T5Xe9hzdzApBaUHF8xcQIqnaX7ivoux95JK69EdKVWyDeVdJHQFkNxmnajGSAe8URthwe/6vfYR
dA99tmQJWn/K9zhu1g6QmjbRZZVTkhM8MZTltBshjkZP7l9GLcGwTPy6TKxEyj3Ga/Ae9jBwIIpR
BDNWdne21rvJAiE4a2Id4yOsZX1CUdQeYk9LlBaF6xeWPFQEk8y3vZsQE7AigKDzBMh3TD7wyNRD
sW3QtM2EPZPRQF+URx7PZYTK9WVeZAmNzvN9Io8XZhUdCb3RGpLA6jdAdIjZnQecJHW4xvZ9BuQ6
KkCn0QpIxJERfYmtxVLsbKsXVSwIWgNVLPqVrXXSwcyWfVsejUHQ98zqnTAjJ6E5LrBvtMv5N5Ky
ZrQmMyiAo2+0hHam7fpu8572gApoyH18Anvi0DTFF9IZG5Y+pKre/L6toGxO/zoQBaZ1RRaPH00K
v5DAdyoeSwORVCtcqhlELacvTSVLfBMYQbqj4yb7uSTZHl87J8O3/UjhEE3ztNsPIw6B6ExJazUN
EB1a+x00GvpiNiuohDSukRl3eTxi+ThjxfpH/F+wjQ6IXTl1OjvyITiK0hMZsF94k/CTC6Cf91ej
7B22t2KOcGS2CZ6E1q3To26S4knlVEPaXPWBlzNNV3+wnpuPVALpj6PnW2F0J8gtxzaELYIMzw+/
sjLMjhI/rHDhSfIU0ExqJDZr1CYHdGxAW2BZDn4vxrm6BQhRV+EUTqVrJ6MIWbOQYrMG0hKUeXff
9/wq78+eZl8yY/sMPfCBpgxOXdOm40rFLNhuNYwqWwoRq514kkkP6NeSO7nZMAC/B4NS8cZGX5Bo
VIbFxIYRAx+YcXRtNT2JOZwREULXjZXD0N7FA+dGXFUBTTafjBSFNNXcI9QOa+wjW7ePMVYT2HTE
ElrzQudn7JywQlByyrTUbPkgs64XjD9bZ5G8TyKmX5wRxjkKsTrtIHhbJY+BbFinTvKU3SPe8ojg
kX8esmYmjM+hhbSBKLgba30AmSyPhpU9ju0MfH12vEHLyB0IMpCexjfRSm/MU7CfVl/F8M6EyEcw
9GOH7FJgzi9qN06uf0pw5GajiX03M2wApwa3YK3kUD76Q5ipCYmiQtzPqEtSrwwSNgw8zMcMWXG4
lh4vv4gyhl2d53Lt9D3GV90JHr988vw/nID848maw7S1jkVEd2HvYBietHS9mzcF+u6STxZ6uubZ
jYVlpCZICXkD2oMBh3ORl1jZQJyCSDZ0+UUT81tp83C1kAx06DjyOVxrN62X/UCQmikOymrvzpK4
al1iZc/snrSXujf7O4W7RTOMNAYVQ3wQypHcVBDsj6QV24HilMIjvCLdoCbVhM7YPdq9HR+51YAV
3By96qdwq9hnfKH++d518d5LZ46T4bvK3+vgELZSxuxvEOZv1MNBPghgF2fnSs2it7iQ6moSQLWP
2AFghpMZ6iqoNt+8yYjFa4Mjk7rd90AAEu+gyBXflkI6KIR7atxJx/9fC0wG1B9kitHQNh1JYoAu
J7BabEzVUKGKv0P2Tg/6IflTwodhxs0HGXrNqkKR52JBYliKieQy/VCG5etFi4PRkgJ/5scqsyVX
LZ8NrXVhGwjrteb75C0yyWHe4D1R1XpRbi+V7S0Ysnh6JuGng6ch95Kkg3VBRh0tlxg5Us1RVuib
+qPHr7l21qfhZ0pDFzPB/gt8pmBeqnJOkJPlqG2FiAqCYtyuWqlFQtyXo1UH6ONFaBVoftRdLgGl
evjulvqVt1jIIJrLM3cyqfMNdVz3KYtLGUUI+Jo9TgjlndtKpaLyCPQTy6tnalvsBI9yzV+MPqmE
/CoSXd0i+rKNbXXJBxfXQ7Z6ce+wnfH5S4+lxutdh+jNEbyE5FtJPnQH/hiQ96vtlsw8FnoaoMw4
fpQMFlSNmeUNAtC217DoY6s5F5k/9TvlVip//zHJ16qmd2fjTiJW2n1Kp15xf/U3epZsYLdlJ5mE
Kr0k3npTbTVV3QBStIPu0GFjNoblE6YFHn2raIF0htvtxU0IUniRmV9Uj5bq/+m24q3hkqa+11ZB
LyssTnAhfb4MJQFuA2BM7lgUbaB5p+E4jrC3lSLa3HibYXrmITBXT/AOD599FXmRM8MlAfAXGaOC
DqZx/jll2YXEBMJU+sM8cNTfdRIDMPBLiL+/IndVXRQkFwgCQwZviX0g0+bccJIucFRA7Up8l2Tu
N+hT0isQf9R9N8LLL2PrQLQTJTKJKXg0e2V7Fcu9gbploxFKc5txKDpRXRln0beInImb3GSq2fMP
UTyly0T92Fs2Ht6RIrdjqT+oUytBDKRc4uVNlFNdrEER6tOLHerusU29RXVfQwNfEfQJFowpV1BM
wAyqm/RbYDM6CHTi/wt563TCrOdfB1bcZala+XdAjwEJhEZ/FJPDQGIMtyFVl7UVHUGZurQ6/iqE
nb0CpPvFujvl5ujLKfAvcH2qvDXRwuBCciHyOj5GDrddz9/vvQChPoD0ObX17ixiVBwgfjp9DtKY
IenfTXhOaI8DxeE7Xjq9egSFM0I4q6yinMlosTdAlL+66Ux5YlG0jL71c3KkXftLcJ2Ok24nuwbJ
CAdKD72gSwZXfjZwaBCS/qJ6DeV48FZ14rfF1T4T0nkmv2es28FeavJR9/rkYyfOHQF/w0ZAYnf4
4n5GFNCrFARumGLczC8n6ZH4UmV6oMhbzrLQaOob+/9+seiCetSgUaNSDWJBTkyFoEgxDwvs71Xf
a/+Rd392B03YKQygVI3BYKYxTg6AZrp3wBU9MXpNY5jNCdg1pC7pxWQ6co+wjuSbm4zUd26mSiQp
T8En50V2JhfhcFUVhzaNLKOPK+k78NqI5rETE81S86hsuFueUxDDCb0utZ6+94/SFTVD1SkiWhMw
oGG+5ZhqE1IUSeqFKxfHtPjHTaTqYdEw4ovfm5I2j+33qWNCYlWyCFhcH6g1jSKeDl2M08YaIkgF
VUl/tqa/JylF12KRiMnnMFs/0spnibCt5uHrOZ7V8IQoyHOaRVWSobBUOP/vhTFm6YV7lsGjJS0S
sCQNZq/9oxDkHoYXpuOijYyZixGDmoDboOcpPb0yl/yW5XwcmiV4l4QwfzkdN6K+k03rQ2g5Fnzn
1BTuo3sRACDtb7UqoOJ8przOt6mzJw4Nm+ff8vkTgCgdAtA50Dzey+PVYgMTgrM13dzIgrh3yP2g
3hobZ0SFbauQLiqHGN0XAA9w5HyG5ra23rV6b4FI2LEjhnbEIFa1WvjkzkGIZs5RWU7B7Ay6g0Lf
RDHNIDy+QKg+kg0a7fo3h3wZGDpMtBOQSLOQzc2RfYSk7FTjhyhOaDOJJ7TrI4PvcJah0L3wiDjZ
zUfO94g6EK3hUZaAtEtfrpgSi1QqgWLTdEYSbrKzW2OW23DZiZnkYRlqM7gGxPZAXdoBk8YR4A0g
dtfNrRR4kVFNtDFMo5YC+oasHwniqnTAdq/h0eORN57quqABe7Rrb67xoBqfwDem3mKXD+JuIK/n
FAB0rtkM+SPeNA2aXYQG9b0U62FtK7PQqqDGjRn6a8IeXb7oFeICrZNP1oyaViiDhzWCexh/kfj9
jUiZzTfE9sPs00bNpAjuP3g/9C5252GXNe0Z/lNrpNNPx0BXahaNW1BOuXptLCxN39oAmzLOzhum
YUe5kIBuzyEIXskGl45g9laeUtV/C6rVZ4R7y+2lhsbjvloKGXS0+2ARakIZqXEpQ1DRP3Bus1Z0
Xu3haInXBz75PWcf2CJv+JYJYnJLchPqM7GWwaPzszipE6PYrgDiRaPjYyFZ3xAbMBn9AxmIiDA3
m766CtNMsOfpxuyZYPAjG0HmKpV1DqFAV57S252tCN3uxQbvt7nhY6cKZk8k1Tqstlxudo4CwqVo
K8PVpmAgPPplvuyRcxq2HhEP6Nn6j5vj0PftNbvPadEt4gaxbs42a2a6n2K6b8XLfS9+EP5vjoSU
UX9Zhe+DDVXKtEGlb0JDr6jws8HlOM+QoT60LKcCaNNU0uP0SQ1SFCUOo0g90Wtn0YvK5+gfdQKB
llTZmvxTH2t5uqNTTPgD97C65qAoWh9gA6pxvCVNqw+Vmw6rQMwyvvOw5+HXFGvTD/o7xLIvGMP5
SiR5UPu3gPxSXM4sGZPUf9Zk4Une+zF6qPOwB7QAbdoMc3uHbd1sI8QL2uyiMzkOmQnx2uhV8UYG
or5uxoI4Da0iWqVO/a3CT+k+fFDMtdp+rZcCfZQdkKPAwe9hmLOf/tnYYSP2/ukCYxSsiQ182gp5
lZdqTPoQOxTnCioFT9t+01WpN9FPvPf+/Y1AMVWTHQ7yWajJiVLvlIVOLPemWZsLJtRSPmyuy2QD
jnh2M5p4pKRgjDSwAmPR6eSfnTeuXWLn2ffXvbbF3CrLPX/8u0wasoT3nSomKgV9oGa8iA4/x6nn
8moFGtPhN1L0fQgfXHriuriYkIOxmam6TZMKbwMbkhMT+RoOWn1nnz89bziVZIDEH2F+7QMUM2W9
PmSznT/XjA2tbxWhEIBr68BGLjME/ptvHGVOpIJBj8C1EGvq4FgIdsgCjjkKD2S5DudVm2uQec9v
AJhmGJZdryGcYFm1DB4YqVDWGCB+nVJsC9TCZusZRHW33AWrjYt68Kawr57nadKQN1e+oq0/MPhX
RRty1JmenD05vFTo8XgS7oMPxLp9D3/3psyJlnGXd6iDpNS5Qudi+vzIA33YZJ3ILPLEEeQoV3Gw
wmIScfVwnTdGoFJWGNZu28yvfCoZCc85NDIcl5WSUwekssQCBQYMxmQpXj3SWN+j60mH6EcrqLQK
DHa5SAX8TwugmRtFI5oCpWT/M+BfaFoxoPbBMCf+rTe1uTDaWBlibwpTBE9yA3a7Md/4lTuZwbPZ
ajPsyce/QING/ZAooabs8uDYR7UaPkw3zTE11KUjp7nuH0+2QIoT6uxVWbTXudQZdIwPngKPBAn4
gd0OuGpjLnXX7QZ5OiGw8L8T7AuGcsrPM2GdtrgBJ9yoCTbUslDQCY527tAV+5U3phNQM3JoFiYG
YGqKRHXBIzlFo8QVkwZR/4SPmPWnKNZdk2duxv2cGaJGQd05b90AS3VAQ3BZ9aVfVazDx8DuYwS5
v++nHO3M6/F7vBYKCeYUipt3Ya140P7e/YRo6SnpUbSqKruRdBOcilM6RtVgVaN6qBurAnaGIO9r
QtWfKZAXBVh3RJFEdTf2fIMi2jIb4D9lYut+NFZu4y/6AOnksxWlcpx7r/xyCtFmGPBzDogGsQCT
HFuUwFFGjYy5ce6jRVPYsMIdC6CoISiwHHPLn1j1RvurcHs/UwZLFRrdJqqkDPUjoBN/Re/pA8Ec
Gr6cCracmUgBpCEyR9elS7sfA55yDpA1CMqyQhqQIXoeGBOvAVExDqdTI6/bvhymTkCtdC8y8g+F
VvPmgTMcnnsSJCada+QtxL8Z5EbFnlSQnq0aRSiirHQLmPMzrf6hO73dRYo6u+AY9c54U9+1OPlA
O+x+Gb7uAyYznkc0yZ1OcmG2xxYaNurlRmaBCktVZk3y0lhD4w+IvpTsk41XY9mBALroPOX5MzX0
RVochgq03OMKvgGKN2RIlJnvgu9mfWgQNZ5Ay+tG94kqg5IsflJYS9fCxu0JqICs4f7n5Px74jYP
cUJcWT4tcc3sxk3uuPn9h9UY1pptlqSKjV8BekeaVsPcFXzbigLDpVA/AWoA+LegXk6FnVgO6JRm
mmNC4RkG7nBVazYiZcQGCO+6XkTAdR0zNGD82ILsSxlwWy3nV7N/oMMzHbFNfrAVTs2fnRwixENH
IWwCl3G9ong/5+UEX72UzW56n8QKX24zy9tfd4l19cUDZaV8rxAVXtNy8hdxeHerLGtuEWzdIgoQ
/J47UfEP/mkCZ5rnQeNGnY7nk3DNHaBiKhqpCPTjaayC/BN0yFseZm7bg91vm+Gmuyczqq4xBOdr
7M+hZK0QWq60XrjUeUnC5pfGWL4XO3AMd7+HhL485G7Bs6gfn6xMZRfJzgsbzpyUQa4ojqG+P5d7
u9gbXQuWcjq6WtDnk8TV+kiT12P4ub/Gi/IR1beDMII5+dk4OJK3LW6R2KzT/RJ6rEaCyLiDcrjg
YZfnIeMwCDbe1sJM1/EKAyB2RvqwTEllr8HXMGrDO7kzinteUaj8MkuO8ecmbV3SitIlEUNdaEZb
9AaMHvf/K2yNslZPYVzLkFJdlclyFDbTW3E7I/F1ryNTOH+QNZJccwRs+sbIyF02AP2guYJepkHx
JfanY2Mt/8EC+uZysU5eUNs5cGpA6o50SVTvaPp9ZzpGKNaKVOlnLVI3o7+eBXD8t6wPIrfI7hYh
Jng9xQUJSCP4RFTNH5ykKfG2eoZT6BNzmxR9S65xGcoGhauJcf3S9T5GIOl7DZOTfv2nLRMwaWZP
Y73qDMu3JN4QHj505S27M6JQbNnMVUIQL1gMw/lf8vgUfnEcKEIe9ZyATXsfBoj7PmfsgFVEoyH1
Zp9g4anGKM8XFrss5NOhu2viwovf7+Iugc2lRamdRRSlxVyYsnqP/x09856g2SG8JIxVOb/pmAV7
Q/I/lHT1Wnttf7SNy8C+A5Z86IBd5dOZ/ySMNoltdCc4gsMAHj3xNp082n/XgEo1k/zyuguDUfN1
qUmjG0jwjl36a+KWitZewsOptrozIpr+fV4MD6Y/BK6PpoXR7lfS1X2C/z/mwf0nB5MqHAATS7zS
YMW/trzO+oqqekZjpZ/manyyn360vW4Pa39AiApqfqZRliE8LesEpZGSLeyagpL0QRj1F2Wxaq8+
+zc1rPHUpGFqJ0JPxAM+26/mpIxjsgrI87k7uN6/yNQPpsDKNWm7638T6VbmOK4VVFw6bCHCaPH7
kmhrpftK2laVsnpLMdiqFqxfPGl1uL0joDzF5vPGDNH5tdGg+GEqlSGO8OXj0EfOnFjqa7gl/F/d
7XdjiGJ1CXwvpIdDKrlw33c3Q8iUBQMKZUEskmRBLhBaW7IFnlQLwXMpQApnX9O1RAQe6bYqkTuG
2hzBarTLaZSYvB/EwTWeAoQXlZV0uTQ6b99K2dFm3wKIxAsKsTmOj4gHiS/C3Q+rsQOQ/r8UUT9S
toej65pr+ooDkh9aVfWfSL9MsjqAWwcyIjTsPcmZLKI2gmcj9SvAM6Y6ySO6cHV+NCKnM71VagoW
3pGwwcGBYeqe/38On7+/umiLnYBrSjz/TV67X/LhNES/YwSvJqXbQiCW+4bAnP762u7KfmKlM5ZB
Rn79wIg1ZTjGUPqXOfO7cd9V7mwY8piSbrj7eUXr97NqAtaeZH7AqXDB4MuUW7cQJIloPHWWFxom
iTsFafAehZM6JDD1I0qFR6em+7Y1BPr3y3o0POpTE1SgILWN+ROI+gtROC1FVksSGO4W3UAUoHFS
CkhPVKp9NUR7LNs6WS10YOmd5XiZdEq2zhk+z7WtF4AX8OpurkpefGWdXvstIFV6SwfHxYiJgUiO
ZY5aoIvFSn/ZpBReXPayuHFO60wh5Yg4Fpe2NhBIMG46vhTM12ziLLwOqcz2sAILI56OgViushfp
0AZOKl2pz4e5s02QLRqhV2cxnKPhJD2R2k0T2WUawDyLV7cN/XiF/DT2DGlHNkEFH7hYQgORk0J3
Gx4Z6pCwH11ealCR1BMq15F84S4cZXxZmfiEIEHPbOz0L1CcTO+/Ut+yKfilRwCKJuZbD8FDJYgD
PeExtH/CV4DwPtlXTL2NtqkG0UsoPwSQopZP4CFZ5WftPSx2N113gIaUbmcgpoTOlsICKzRIniE7
ZF0NIng5Wat6XU5Lo2Pr0rEpk+WVBwXc3kRg0iBKHsQiqFhS0ZqH5vcA2J535dAQ6gEhBW05svpb
XtHHc19dKHe+ziXg7O259+IEy+lc3P32rXN2FaJpHqw9ZM8BIGPTlmkt0j8sXei/X50RP+EHyIob
kU55lMTre0ohhW0Xe184Cl737/w5G1iUcuFlGVVg+nEtQ77gYqKjIt+VCQmaByFPWSoMeArHxZ+o
baAh2ydn8Gmwfi3xpI6/y75EJQr+g1pKuxDxlj3D2hnhsRl7lWQYMX6QwK9JQb0ap6bNTCs6Hqg+
xO84BpQXpVD+GZ+lgnVG3Fx+sk3+z2719nRP5WXKfy4idbINMdQDNFVrbwiRJNNIT3/MHTJ2YdyR
RtZIyf5VxLNA/BgiIi6GBEXZz89spnUWrufkwrcls2Atoyn01SEraSMhiRdhz/dW3mu9WyZdutNz
yQnXKwqA8inBLjnKK3DxsCJQfkul35NvCrqOfQaXBACDxtiBF0bi5Yp6VHIcptixAra5ohldtxCf
TvwLA4W5CXca9EX6uG3MVCMPU2wxHhK7EPrUlcnEQoCTnA6DFizpBKmrnPlWeEkSjeiLlbXjMgRb
bU+PiJrvDENCR1sr8jwkUJ9MLnvi0MxsgBbfOL9f3wvvb7J2vbW0HBBnoQKncpDLgn72zFyu432Q
spJuhiy/pMoQNpU8X+s4im3vz/xkmJXvHwJR9CL5In/VCzRKkT02OTZb1uZVwweuIf4/aI1MpUtz
9WMiSrNd+SaohatJq8VDb34GxvQQN+xBpTjhjRjLe175wNLDOV8J5bTgaRTgtU98MJlxXWT9iUXx
Udyv9Ans0lFI/adrycfsknI8195N6IfKnmXxFwNhRG0tJ0J8taZVHQB/Yzcl6bD1K/gjG5KudVSM
p/eKwdt/3KMOqCF+GW6SrUuIfiIqFkSyHP7zb6L80w+g9wcwiJCLJn0CoQTGIXbSw9+UNDdlowL9
Ih6XAYY+YVYIllWDi/YQ3Z6mzbqA/0nloOjuH9i4P1XSJFFK29zCQi9XxOz1ll8h3dAR7P25mjuO
59rhEA7VChyWEn0akkjgKfB5un0mSBFTOEyZHsEkaDP8XvDo/rMoJcqubI/xUV1o7Ail9UC9tFcF
6idD+kOVMVtl0RjFTiY2AAtIbArH/XEpKFPF8tuV0RQ1ok1mFDRvT1UkV4XKb2toiCn9q+qfv76w
EaheBOqCcnEvr7RSsfWPUQjaT78gonNzTAqrqp1GOuuDjRD/jBeH/wVVvF9KJa64ymIZYlvR2kSM
lgRlzklYz36iDcHC492SV0yhQfnEwgz7vZTyvvMBx5CvX1xI77f7rWVjxEkHXnYJerCpZmopmu98
afkRHGNKrbV+ajWs1bK861BbXGm2z8ZYWTQa/7wk98MS6jfhi7+WfDKxU9iX0ejdDLe4oknjc9nC
NtMP7MZhglQXRpyJzs/cfYg/G7NayjkFua9ahB3VBWJUH4lgC3EWI4fupHouSzFD+I6KQni4tWYB
qVYObW0qbn76T/SD4EvVI4/AgomLVwDjQqpkmc4QWMDqS04uSIepLNGe6qvPtmoXRiNMLAuhfBgZ
h/sXTtOedSwH6SX/QlUUkVXE3uEIqN3bsKyfFj7/0prSn0V5cORvPynW38/O9ZlMVwGIYvEatcwn
ZziwVqAf5diGmDvbjjnBjLcG1UXFAWami99DzBq+aCgSm/7DdWaKoT75uOHWcDcpgdV67RljHaVv
RLjHmMF7FfaGg/8II3asby9QdbXB2lYCrnmpwukDAT3l9UwqfJPr6kTj725kTnNV+u1ZDWxBqfHV
0DMgP6RrlsN7XF2r7tUHtvNCtMdcwRcUjbRJDeOSSWa4M4YcJ8Jjln8ydsoSar+QL4BNRvtX6uUb
ARO02/+gBEAZhPklzIvA7E9IZDBvALch72CiX5Gz3D7To13N2GwH+RT65RUf2nfoEtzpq5CQVyqx
18sUlodt1VOE42DWc++dwEkUs78WESIOVsAHBEVRiiY3kFvkvcvhAANUoJ6yV8EpBSibsY6WykfZ
YldNH20vhAn7ScJASLYHaxG+dOfbMtCPRbF8rlwUi47YlXRyD/CmIM0LLpKkvfy2gYKLxQWhmF0/
tknkG5hP/te2TWhxsGhlB0+mKeBSFr8sfVnfmcr2OdsdP82+dalAimjoojfsqcV/yeOvxxd6vUtB
QKgTzSQOF1xUO4NrA3m44g6G1T7CiuI5dZZi9m2i2NxEdm4MSKfBBmEhLHbbBslTdiXTfkVDKJsx
1oJfH8A8/tUByERj6ehPCjHUw1meREaOn7w9ltacS556pEJbsLmTrdkby01D6SGlIG4/axh/vEgQ
j0neFwzYgzYhTea4F0q8W5dCQsMi9/1DBsbaTuGkdYnNiKdjycW9kT9FPjjEiG5GCAtzwTllfRr9
bpXb/8HvguZtNW0sU4cW7Z57z+5Lmmke2lR5EPyUwMDhCfg2eqsPsl6gXSPlrKCG5jy1z0py6nDu
bVuEKjdld+XpmvSF8dvZy5VW8lJ9jMZkq+4JJQWvzYUuzo47Fkz6//Ou31Yi6HHU+Y6xJVex+l6B
0MfP8SdtWg6x28Hwf8MXySr1fP6G8T5frwEyOZ4XsMEHpjHlryp0k3KNjEwCkZLRA+la3TJFKxUd
QSPKBJQ8ppcgSNQjsM2QwDBXs3ZidlChv7RDIViIuK5Kt/huTj2GdCQPzvFCfwC3lZfetYRhrPph
QEZwaK+3vIRy7kXN7CQOO+QO8J5pprVbz9U0wH9rgrUTRSJOSDNYlZVtP1zhgoNrQ8Oyupo/eDA6
Lt3EiPg8cdUVkWPbUH2xImqoYf6qHghLEYhNpkAbTjLsBNGnxfcNa+vRnEthHIQEksFp1q1gv6e1
fdxgqFNYQkrxjEgT1GS1kLW+KGOQBYTOTs7UMML9IKJpbof7MNc8O7I8ThSSW71KQFMa9MT1k63Z
tu+VVDLgpdKCH9wYNPUuT7B0rAocv8j86U0ukbE/InmuCsDtkXD3UqHGJAdQpELCyLwmDhv958Rv
dAZtcxdRFJd24s4oahcOHPVqOhy+80XaYHRaLEtaCuCMfzyPV2ArexiwZRGox77iQcrhI9BOnbvM
MD8ym14Et63wFe4SFMCDwNS3tbYjYWGwt+V3WacOC5ffK0Pr48fLBc6fhDK/FL1Lz8xuQyTDhoEO
cVCVRUtCPgMHycXiWkuoNOIQhQ4kol4+i1dBPjAc4Kfesx7Fbci/09CW4QHhgdYu4531j0ihlIps
UIipIYLQmncWvM3JzoSBWD+a52d/i6Cb3lP1mAMOl+MzU9Q5Tk3/8fS++jGbJNgIV7hrxT9e07Tr
itD567wWNXgFM5XJg95bq+yRFyK4uIGwDfLsqJKw6ywLX5rOWfC4ZhfaLeE4n9H9TySRTVpKLRFh
9Bt211e3SdOjKT+swKXchjKc8Rbk2YpIGDU9uYeTYzE6Z2fDR8hidamS9/gqdkPWi/egh3ouLyOT
KJNDPR1t7BMjJkgIiLKdZGr34AN6ov+kJEKYMjCGaurqeHdbTp1F0sEyhQ0nKzVKLPz/YKVw9Oha
BS5kT7OSfpjbf99dRF7Cmr7c19LaT+AXHA8CU6Uj/RZc+CIFMf86ojSqdZELXVSp2z65imMq+GbY
NYsPbwi6U38yxMCNDyZRBIVpL3Puv1QhJpFwjsfn9xyCopfcMl5P9DuLWtE7noRAR2jbWmsKtS1x
CycE2DnjAsiWy1zUWlEuwj+Azi5wQ46+zOe2RPkkTa/bm0gJ2kUyJPSDGVO7vEE9woP0wP3TTVfy
MoZM3oHVHI5onJl8EsWHYJGFvBJhhr4jmhfZ6bo/3tigH9jwnDSIJr1i/jo5e6aDgSARdUTVgO65
FnAowLiDTQ0zISzqnxvq43CJ1y8eTfKlDfefoyvBITzXM+zvflCYLHAGCsVf/YzLarGW44zvX7Gw
d+dDsGv3MRrdnCPTg89y5iH24QTtAHfyyGwK5f+SYcCn9Php7xRduHD57vfyziiVkWFWz8NaYQfk
v2ybxjEaOl0JiSCyveD4dJcMpmu/Ah2LSsYraIJbYK1PhetMJA01Tuy6BTPWagp1fJNUaIlb7n5Q
eVv/QpuzK+1y8AYP3n3h8aPq6mp4n3yN4uAEoACNBKh/HnwBsdfeKU9VaHiYAz03Ljg38TE/oEjX
nlrZ37XaeLgMX9lg6lPN24Br2p5grx/kfqcP865fmFblrqGexHWt3FwtOfiIFlioMDztIH+Y4drM
O0tW04sJ1mihWQuMT7B9RrRXee1XWjjkSjwjFYvGoELCGoeP1R3mGJY9rH4AK6+zT/LHjblPcN31
xietczIE/Wad5fTh9tUbahFtgsEqP5rsteVr4ia+1u+r6B8wFYea9HjGFK9fNDvGBbbsOLv3oOrF
HaabW+/WmEWvXFuW0vUFRJxndcK3fI2Qqc2jW++m0MJ0q1HOo8FU7KYYLDbsl6jTXq8k/g7nzvwa
ukqP/tJTS7HSqf6HDvjkElCgu6jBL+GuFF6LIYbj8URZCDAusPgWYFODxkfdZpMMLFHnRWfDZ15+
yKquqvYfOEIavqRqjwVpOb+Ba96oukEI1jad+NLSc8nPGlJQKvgFx7bkMuRQp0SpbW5smyJYYjeQ
Gkb4TofqnJ3Ftqo8oAgYaw5v6vaEXoTfREEL5Hd+jyMTa+AuFCRaXT+MSINKqKasz0NntVZhQlEI
cQmWYHIESIPSshuaePR3rxoR8DCoYmAmG9epSHFEWAyeEbJSkRqcIT5vRP/Z5bN6z/irtYv6278F
cgQ0OjvVFk12l3a26NfoYdNPOyVXNyF46c8Yu/fMyvANJ8FIm9Es9dMP4UfpsvuBzKT+r16L69Nc
by37q27cMGhCM91e3OZu4r5x48xhpvergiN+PvUOsn6o4YWWAObbZilsTzeV0AIUPXBhPeGXIpil
HFnyylpkF0VACqU8zuhxke+kWh3fxAGFgSjA91EzgdqZ1KezHhKeW+Kwso+BSbP1b6MAmujCpeza
441wT1Z2PaaLySBJHhJ3TAsPOYcdEp2GezH/ca6btigJzFHDVeP8aKu/7XX0ublDJ8RhEeaXmPpG
U5v0VcxBIJVwLYyBT5Wy+AzRXXBTt8YUXwixRY3/0zzFvW9YcD46CtzLARF9ZfAjnkNu70LU5qV3
wUsXsa8rV8eBlmCZsxoHkzMgr7BR8bJScuLvetEkFVEyUdafOrkCXfZk3L7j8L8Mae127Vd6Xab5
FqhKQKnMwDgdrHiCz/nAhjK0/h5jVNZkDgYi+2xXtDDGP1tNencCThIHiFlJayEXQq4o/K79/2zh
NzISBMAvl46d14N+NiIicdU/zpUuDJZ13fbnn34MjhOIHKWz8HYwvrr7BJ27YBrvyFlKJWD9oDhQ
pXwe91Xetda8qCAonN9yIqnvytVbhNXLCw1Y87rRp5QnK1+EetlbUzRGgGEsLNM3wxWuMzpYtT8z
c7CydFXfso99WPV40yxSoHcTvEwaHRl6B5lZQ8YPuBYlbGjOhzJ2cLf91CI7x2aauJ7MOTJSQCUL
LdPYWtuqGugIc9E48ddTrJspuleswyOjaL2mnmPnhlFRunq8cjhws9kv+lWIGDVh9QhgNWyAa3Xh
XBV3ahw0x3dro0spHToHSpham6FFlwtw0ZJ+LwHomIbX/2vC01VV7sOCh70o5DUW0f+C6Fi2n3o/
+wWaKHJw2FF739QsoIXUfduBAzWObXus6ygdV7YUjgGybIf+BsqkQxfjjujzE4S78T7TrMg1bShp
B8QQaJ+gIOl7ErH1GPGdz79gEoZs2nOjYhRh3AKlo3BTx2HH4BnnNDLcNRyqA3wn7Yn4trsHKpDT
ELKQPdPEOMZXQYiIVmor4zawoofkl+9wBWij+ogpquyrSavC9l4kMgNVHAnYZqkCumbRVKykQfyz
a0M3JbAeDGyani6GFDS1zp8rUjWJoODbayiyZZaTeALCDqEtjhLhJZ5FizBM1ObtvbH+ez1DQ6XS
qYEnoJU7qkPykYll5U82JsOj3L92/lKJ/mULr8DxTXL9Om9RiFZIU9if4gBmsMT7vfdsLnf4H7D4
Jh0igAAGDmmuAGsRFYRCIyj4t0JjhP98gTQ9r28nd+d25N0IKrvdpGFqtV4ApFBUR+STlU0pd+bE
R0inn3oeIWxX1Cy9j97mu9hYbo+Wu0If2RAOo7nEJsqyFKZkP8enj7D5ifxoXQXC3e3Pg7cFq1JK
TuKivfDdoXgMFeQWJLdujuR4StiHyNorTXrkeS3p/5Hc44Tqdm0fC2/WmUwRRYftmIgygp8NzUej
ahm1j5NXxrXtu++d6PjjycOPEZ40wE5cgFLl8kRKq0cpoy+WFEqZYTp4O0/qbT6Lr5UDW1/CqyRF
Ps0AhmvSpUHFLEp+/MP4cn4Qd5B+xPh2vIy14jjq8O3hZqpj0tuBakdXZFrGi5qVP5EkVtLlwNVf
kqewn3iWOZUX7dtwvInfrK6et5/7g38ASRJvdpUw1JoDBv51qSMxYN7OpnijpqhyjB3Xh1VECqmJ
Azq00L25VAmUEUh+k2NZxZZSQxO4fWjH+7JylbxgxLQSmwCTgVvIZbhWH7qUXKq3hq+UT6rkBF53
3OfkOO7dni0gDh55cAW6QcBvjIbeTwc1Oe6AmfxIRPSKeupg/vrj9/DwU1C5LunbnLgfhkgmWn70
+kPnRJVCA+kYBWdpEzNEL/edCDl0Ab2ZqZD86R4qmL3xH/sOjesbC9z5pKFoWaN4qjPI7wJov7fn
d5vYSkTXU2znBr2VVrdSQKm0gGncn9KEZWO7YPd9ELdUu2OlUm8k0E63a+zWV/UHWNj+sXpOU2Ok
4fTZhot7JfbGuAHQsLJVGp6YOHWxDbvm0mw8YnZ9X+Q8dRbsLx9YwLdkuWh3woz/0YEF/hf0wdQD
zQEuB/rWJJVI9RGQIj1q791eNFKZylN59LGutuKE+/NHQUg9jnQd6WxzbRbi7LJfiJcoadHlAHA9
SCHUQR5fRam7hYydzWf8WFb8dx3TlSAqd3/klVE0IAhytBoZ/eN/U2S5xgsamz9JCx6k1wbuaA4k
y8RkZ1E2jmVxcQdcI2qH7RDK3HDfpgSIdnZe62GcoEz/k9IM/Q2bvvjvCoyEfR0+uKlnHVhIK4J8
jJdw/Hf9O8pByFV7KxBKSSAcwB0gkVRgua+UawUO0UnkmMBF/YF95hT6orHzsig//krJumKcvTW/
swazGO3doWD1h4ZvDLrARgVqXCUb1czE5X0zHRg8QB/tpMpCf0gq/wRLQVoAvyKo5EwCQvWYaHr0
hWYNqhSSGW3eIylVwlUiH+FQtOcjc4vNIT1OX+6Pc6j03ja0SnI6ziITUJBIj2ZWYw20bBKZSPtE
1zRgr5v5z/axdpU+neCri90473rZUsoatBgZnvjLs4jPE6Er4p0HlOkkVaxCYiVLun59/c8BTH70
khhvfRSYKTG2tsZhlM37lPr8BRbJjxpsr7IE0lgv3jtWbqDEd3aFiK7WOODCOrqTxmzfEiUIoUpW
K1TwikYbW7jy5kfOv9JNFOztfXnSa5LJ2KNY58o2WrS3NWVq0o2RPvUael5gblwLkEC/KistATQ8
yJLPnP8AjzTI0AxlnZtCe11Bn4jPjIFn3KZ3cB/cN3GsD6jh79lMNVM6aiZd5Fv2DBxmFhXidAT8
HKxzc+XyMFDra+tvj/UjtVk19uBw59R/LtPxTDu/JjeI2of5JIiz/8N3uqgbjjvc7bzqfFat+aMx
PWr6O/KEnc/egFQu86DTTg524EopsEdZS1wSxVfYwNrRQT9cI60l7BYENYcPqBLE2vnAxIrGDPE3
xh5RfIyFUTEGLvP0pBz5c2FTgWyNmJEhnlIy9SihE49fRyZVRzhyZBKmxrrxcJdZgdC1W6u1w9eF
VNpi/FMuIDll2x7Z40bcCla/RIGy69InytH5NQH/KnHIUU9Ev6i4o9BZho8ymQyfvD11xslgxUku
kd6BePT897l5uXTTAeG/t9C0U5dk33dlLscQgsNxaBqjZLkGCZ18aLygRDywBpAdfjSQ20DS739P
0QUoBtlxuh6YP+yNc/1/Ku/v0JhXABzUdB6ZHJuJnn9ycckRHZuI1Sh0GaskLHRxDF1qi4xAfT34
J6tvkX+qcTr+Kk4nrx2htMwsJYTbbx/V04XZ4+bdXZ8h5TwvMfkz77VU+4ubrXu45utGURWR/M3G
LIy66nVEVZS/qdRVLB7FnsK4w3TojeVnDz5EZG3ryLgVvEh3aGP2hFrenzCyLNub1Tfac9+vH9NK
s3TkEFcCoB/ofCg8BYSYrqirgo39L4brDJ92ScXvMi6YUWr8fwDJ2lUtNBioqW+LHcIAhgVRW2TU
D9kZbqMJ1j9U5NdMTJedXePH4465ILmQmleDBA8NH+QI1U8mgZLL8aMxbHH2TOZq4SjhzXeF7tzd
Q+fzUORxsOAUbyC41NcW57qBvXsIT9RDKqa78fWua7J2EOpN1WhF38bG4AxIgm8RLCCLFtAMQ5qP
PwgMQnuaGSxtoFXLRJEQeIgVVWSZZfNgjvY8YBtpPRZEbht386+TyUBLYqvPX0CxOh+rzMbb9n+k
ylkj1Rt7/MO/8ZHmeYP7rG6Exr+jclj6PokCceXHyA9b4s4fwp7zKXOv28nE6gfDEt94M5fba5SL
3yXxM1t/IGF2DxJ8AIjlN8Py5laOVuZiWtxuuyStwfDzDhi0l5a6yUqtuaDQdHDbpJt67afNqjt1
goj6OU2CcT6NvOp/6YLRDpQM37dE9grzAC0qKZ5lf6VMnUtr0lS1ZMkeUGypVbbieFE0w3JvAvI0
Cqx197x1ZdwP55cpiZVbFtU0iwg/nzbvRdLIUlS7RYUpE03I6y4w148I+S3siY2qDs3foUeGxK7G
N38LL0PGmqtsyPvMhmW4Oya8e3AWYofL0Ayy1VMmepaGrZ9mAUy84nxW4OXPyqGvPDDWc0s3Vg3J
gzxvuA7TbhG7Tl38jLAOvFSfVDF/jlNFWamAQ3+a2cieQHxiC6avB7HIwcTNd8+tjuNrGy7OQzR8
z4J12mSG7UXuC4eFz0ypQkaDjIc8I6VE09/LusdoRcT+Dk6YJdHtjRIgyyIVwBgznqEqpiE4Jh82
1TOeO5PwItuD+mGG8+ccNIYfUdzkjkHDRFWfgMik2NbTrS2E9XJurIGDjddNgduVY7IQ1/AnBijo
OSJn79jnrN7LX09j7EGxUBlc/JRqJrxjN0/NSzObRdd/vS7BL2QtYaV3EM7G1T3ZtIC4YjAs2c7h
1DEVzk4WQGhjLTEvI9vbPYqlvpSRuxcQHzrhV6MP9P58jbSImkeUdfzbfEwcvh7OGwUtcqXHzrka
m9d9hQDrKWzBhBfyv3+H62wpy1ZxW3SHp+Q48RfmBJQk94Kr/QwFJUqQi1/iDv6NDrTJCidqrKoc
ZOY5Etkb/IwW6qTI7f7tXhRXcO/OLNvQXJbfZ59p6g6kdCJhYzTC+uQad2czCq49cOw2eq9OGCz9
TQmmTUdXIPi8rwbCGmcXOVeeVHcVkRTiQZBbzv8n5wGU090nV43jHSwg2wUme2IGCnkTLqGkDoRX
Fq0AlL4WxemGZNx731Y4LZKby1lD0BPj9KAJ8j548RKJ+uC1OpQ2LXYuN6bIxUD4xLrqeIWsXmUu
HX1CGVvKkZeqAp72y3Yigxq0UnADm3m1nozwqukQTPKjEfrOAPYcFtDGX9uIuLfbBqJ2D3+Au0/G
EC194cEA9hxk6+7joYS0Datna+N+RrgqY5KfCU4FEvCuEAxIQtdX60wB1i6rIItcHZ3CsXmtCtHs
TtFiJES6P4RXDaHVz0jQ7OOA6mNynoaSFeponzNODSgtd2d/qsHOuV8JgzgXAs/YuK+DbqtxOfS8
ZyWhE7i7GkXDMgDdMal2o3cCSrkpf4XFH1SKwkjvj/CBo+iITxWa/1yZVesKrMY8a57t3wES6vzJ
YITVAqobR5Ze0YRU2OJE1mR1V9TyK25QH26HpWS91+OUNWGFPJHEGFN41Som6djsYoOZV2FPBM9L
AFOjwoqk3mwLd6bccd8uxnudx5omMQhjXwTk7XVaxXQxSfdhRNFOquM1UXqapa9bRSSQnPBdyXNH
KCGWuTyS8Y1qFyLUGVwTjakgiMqir5/q4B9HYlxkDBigf3srkkWOE3y4VX3mNhqhjRpkpEjPjeOn
YhOi/Z5znY0MyEbREogprlLLcKNQCRIZOCoFhHFWZIJdLTzINIelCwUzxRKm632GgD+UYV4idwEN
ru73rP1GzgcBjQq9Ho1jkQcjxfiJHGPCY2xgoiUp7gy9LU4EAPILiULUibsrjKAYjSd8Wk8XSs2e
Zvf0A306/tVOacMqW1tiWLuZ6ojpjCGC21OVADPvoj34ULLHYBiclNCzFBiH2WIBpsTjVWDLK2vy
VKebiib2koIUin430u0cCSihdTNEXxf8bY8cZtCztAt4KahUtn3r94zL0xPiYu8O2HNyghCEKe6Z
OTVEz/MCYMGvtEwFlXp2PuIGz90eOzEQYHdBnnbyyuVhv0ASyD8IN4bRBXnFUd1+FPzmj+SImZ5G
W3+qjIbgeK2N5HM6fA2czo6lZquoSk3tn8ZNJkDSOosVulxSmAZPUhA3E7SpjMOusTyFo2ZmvJOs
2irLL6YLhEswqLBG3IiaEP0X8SyJ7Rj8AXGt2iVZLYdYPmau1iajYCxkPqPpNU491eClPI/GXwRk
WXLg04R4bJRIPRCG6g5f2lp5Hnlie12mY9gzHh11xwkQlbWEkLupRquYO9eXCCvxzp3TuepkU9TW
Ky9M2WpMuPdj51u+UJwOy/Efyf5VFxPKaIvfCHDu/fJO5fXAaWNJwmn/+3YwIoBSHvuU/BMI/kUn
abq2hxWF3wz/QVM6pmWSV6N8TUwbI+emzkIIu8pFQFcOpoGmvLPrxHTZpYQ61SnJOnpHU+PRuMao
TtjDlpgp9nWQizw6uiSlEdkG38PO2IrgwQlO8akLrdBT8waelZfydXnLrTI4Kt9hqCb18/DlbzsE
JwgIDYAGOrKiY5JIYeu5yNDEH+W1OP/ajvMeMSzRG1YyQ0yNjfXnDVkdFDFVOadnTcTYMkcm0ZDb
ucQDlsiUIZQ0o5yvDx2vJVGQwifefskpshhpIrGCy+5iaWy8JwA5jW+Rahvp/YH1MgCbWUZxr0gE
+Ml+TQgwTJTzroHwGbJNW2iZyUtDki6g1Nyw6kc0zP7viBVzo+LBt4qeeJ5hDAg0PQcqaab9ie5b
LJNSbUS9pTry+XGDc+iVV078htkoOVjKBQtcKiKp5Y4sdcdMEaBDFqVZY9yKpyDkpwTbCh32q1mn
Q3dSvDVrC+5CqlVnj1PUCldm/zFH+3FWadfF+8MtwwPc+hRRJs/5bg/MrUJ8g42caRa7dd4wuy8y
sOfybQj1U99LqdYZR0KpkNRwjf5xqAWlzbnGXPJ/w94Tn1qPuDcq2YS0YSzTSse4E01yHPzeZycY
ZDDskWgoFh5Fq33esGgh5AU9m5kVaCrCoI9mORpcS7yJCdSKN3PHZ+dstClAi3OxpKSDU7su+4ne
8bKJtz48e5eIke26AhDOvMHWcyEkp3JWgM5A4HRCNYJcfeghO8dgPm9hOpWd24r+7QAHT29rN9Cx
M/x/BdF98SOgducS98agQcEeHvSLRGBXDhUxMSGMBNNruklxfxTDYvYUjOmX+DY03OSJ8+Zqk0Sm
66NAPD22jv1VmOF796d3fU4ozVcE3alxJbbvBirffown6m+gNplUUVQBKg+lfFQhGZHaB7Al+Iw0
GVBtqLFMMzPv2I8a2lhrTyatm3hAXw34jaweRnggBo7CK0x2stFjESgF7QrNAGndJsVAhdxn3hCW
bvmOMCNYwTL/OPLdRctSddd60X13rJJlC4DFGtVGqpU/S4eHLR2AFn00aABtftB0LdcvsXA4deXK
4V8wMrLH6FU357b6Z38oJQ57mT3Qs23U0+lNQFe/L4c1aQQ6Qv6LkRB923zPavxuKPmzMk/xlF4C
tSxSgSPxennFBpt4OpPI1NyFNBhugs89j6MIvMbTuBYHh28e55q5729gv1Ga+L9DfgvIqlIBLyER
F02Tx+PAZpn2BUyk8NStFCO7fYvY4RWejbRRAOK438J0rpOB9FkCZMZjv3fs1wvm7Jx3JvLt2Ulp
SzmWUQNz0Nc6jJOum4WpX302+KnVhEqjREXJhT5K1Ozm3x9zqmeXwacSPp3cdn7IX3EGIdLVibgJ
rh2qwwyjhtK6OaIJ970meUYxw3y7F+JLMqTUQYWCtswe7ALeziryn9jIp0WvMh9ryyn3XhLP2N3c
T1Yuqbpt1qDd/JfyLNFQdVes63yGvRwB+/wCzlF9eMKv3BC4TOTponE1LzVk5D57uMyIe2/0NMcs
lO/KP2N+nkhGuvLD7crUHfo+zibiNWHyyndMGdF6sv83DNPE3VKI7p+9SBCydpWHUQx+Vjn07sY4
sxQI6JnvmIBLUYPJe44xQyxtdy6qZ4liok6S5e9OMpkCGcBbUfUTLHYE6VYXUZQcTs8CcxoexmWQ
0CVoQE7L49wXeZ3YG5xYdQ298+qfnOwL0r9gzNMQgGC3rRsBJVWnBiJ9FUrj3lFS0IVOf9d4r22l
BqsR/m46RzcI7KBZjUNj9A7mz7YFZ3/WDfKlHCTIRxTQGNzi+VBvwNXnn/4XQtkbJ55Wh9MUheNT
FVOIJmQmoCeu8RxhBuZFg/riFEFnjO4UEdNCHxhLXH+2883Ck/gnZpgnl+HyPu6Z98K3BJkNAr1W
DYWz6ayru42vF5IY4xeRW05MZII/3po7+wRsuidaPx6MkizopFdFwMPVa2m/xp2V/4KNyROB+wvP
+JhmJjByGIeV+GHpzx5J6bTVCdYXaGQmrbuaUR9za+t6SIQeqXHEOyWQ/kUEoDWFVU1w3Jbs3SRa
PnmQsMJiUpDNsZj9vE8hTDn8AzKf33m1jjJhtQ4UrEs59idch4ZHP/8nnoHJNwQLFcIsxAHrDNY6
YR9/5/XXnN1bg/k32L0qcxtkG0P/Bx5v9GRN4CoEuRiMhm2EGFQlq22HOkOAL2JnNRjGT+NglHk6
UEYDadvU5wiSEg8Jm00nsYX++Dk9mUrrbFzVWun5LK5TE5/KRlVB+qNKvHf0lDS2/wUfjQhUrMbT
BdM5w6SN7mEaLWqpLsX1WNacwFrLn5ypG7Zrzu7Ab3CikfZvzZmxlSxSdNejmqepo0hJdHLX1+Ft
xkel3msOr9DbcRvHFZPFwkHCL1chlUCnp2tvL7he+D4J1KOIY3L2Khb25gK0ENoBUy7P9gdHuXD2
hVFGpn+SXjM0j9+lp0oK1PJkO4K0pE7IMzD08tEmhAGf18J9GVpi4vMO/lca5qMjOoWxlLfF9Vr0
jZghcfHpgizgI4wY3T1YV8t2n4cFhZgI8FCxwwBvgmpQ2jPhatgKrTKFibL7CwZzt/aV/esFPLYf
sfKsskIZsriyIxPyH6AYPP/3FBhoicwH03oG38nPiwGGmrRFOi8xCh3y2W2gm4qMbYWMOFjxVzTi
2JSWXAuDWY3pa1QclXIu2gu/AhJdf3t+t2EsfdzOGcsms2MTv4OaNNhq7BmjCRjlrOF05dRUOyz6
us1qcm/EDjrzHa4PCAMFVelBGcXeWEVe59ONb5Fb3yrH9pmxm0p1OzCi65TMc/88GYTouWklFOGV
CPg11M989S1rgvp3gk6IM0NCoYza9oZsNjfFVj11zU+G0MCC7fH19zzffGmAI1V8L/OV/E7rvMuo
OQbdcc6Kz5cXigFw5isUt4wUFayYBAjKRnWDzTcbFc4kGKJprRUYzA7NW9Cx1pHYrC71pDzXD04g
hyXHTncZmPC6i/FPwqWevxrwHEdAVZnCBImse39GjJKC3Y9wQ97mQtBTgGtlhj1zHMyLcJOnE5VH
II3NNjRpZp9SXmC1hDcDQ1nKAXmMhZa1x+gj+3fyIJfCNwkflZFMrM5VXQrfU3qeCDJWqW5Vn5RS
H0prjHzsjEK5FemDSFLSwnbMi9hzH15Swkw1JQJkR1bnLPjqM3QyYEM0LZnjEYLtCdTwOf6SCzBD
jarS4KpI+LECD2Ki1Y5cD0gboLjeA2xdvflCYWJcgcjGbgHG9G42y3dexW9iqsN+iNhT5XtO3KZL
GtWaFWJxhE2IzkTxg0szc/52dTIw/sFBGpVqA4TM1PSX9QFCFBBcjMZzV9AxfOjwCXwiBhknnyfc
JhNxEirL1iUpD+irwrprWvKHsVn0FBTo15LJjCHWcfgF5i+Erpgw9B+oBf2E1Efd8mklHp4HHdTZ
z8IbFAGTyZwAYxq/anXAaWTAcq1ok//t1BcUI87u3qZv1xDbO7yR0rrjl4ktMJuRnmJkbS7dagig
aBpCF5r/wVmEr6rCcAOL1KF6C5nxXmeTTFukeFIJE2bjRBVk7/MpUw7+bybSoaa4S1xjkai91lTW
j8+Ty9h0nlghMNBgWcGYDTBRLVuetF86Mmz+mMXR8e7X63eacN3wL96bkpZxn1eBGjb4Yt43akh7
DelqkJHJwfaSxUIplLedZQ3VjnHd70bjRhfk0AFIwVUb5qKVs6Au/5mKBfGXnPJKWQqmEEYMgmH6
AEvyZvhK1IX5BppgFXpyHPoDmxOr9KDhbx1h8Sb4RyiI0KTT/LC3E2UKgySCnkO0Iy9bsxJek5L5
XezXMKCHP06U8jPHUngQ3iXxhynFhhR0ZtYzDF0ltOT8ISm0djiim9EvNHKM5LouZmd56sQ2Jd8K
ehLTKab7xn8AIrEPXrcIGrJ4Uv0dNUrjhnD8tg7lKmczJp1fuQUu11qDjfLYqv7/b6OOiE0gVexA
4vXNTDRp3x4LyfME1IAxnxSeQ1OmdVCzvL0CO4y5BPHg+8NLhnZ/J78o/DrHaM+9n3s9q0EK9FDP
/SET9VHEND4MkgJdtFIWpcDIG9ARLTOdqn1L7F30kbsH/Hr9xDr0DILaep+zZchDVtbnUXwQR9oh
S1Vp247pILxcAP+BC4a/ERSmcsm6uLXMM6facK2RpY89tcISj/mObojCoH85q+kctZGshPWHhWqV
si9Yuhn/KczVWoNhJ2kstnZa+x8Kj5J49Xk2d80SQN7FCbtq7t2svuHO4xhZ93ceFzpje1F00X4m
q7NMSQTvLRKnGZeTrEY3cdQv2XfPFeniJYHO9z5v0gQ9K6kOMZoPS1+5d3nRbiI7AiD9aTcPhuaE
oxBe1dg/YL0ZlZKoqyDHFOHeAEy7CVwnY9iNqYVnBLhehuJIqvbvPCaUP7wbfU7xCvneVjl1J2Ak
N0NNPU0AEIO/rVkPWJa4S5TGyujS9QqlAmZxxnt2NSTRLRz6JnETEuKrTph/Vx+QMMoJkea7ExmN
dJi/mkE0u7//vhs5Vfaa/MAe8tzq60MvWMtzLoCV+c5zAxi2WnbbL/yTCRON9rgxJzfdbm4YNkdg
/mER/oy/P+ECN5b8NTM1zfyHzPg8MfGnkl4jZzCozcHVVo701RFRvLCqBHTyeCTrty82eCrGzMZx
gim8XhZOe53JNs/9ds6ndG2K03g1HKCIwrAo8SLAgVc1SJh3NBxk7Yy2deQgaroivu8F9Ed6S0OI
uhpyFVv9VSKY9nrZKCof/vuBeM7+uUKtrH0bCl6b5/J7Qwg4vqWSAVDmZa2BIyz+DZ4D0ssWlzZn
97zVh/+yJE8a9wsnP3DivPWwOBq3KLVQg+PHeBATgx86GT5Vp0krr5JOEQOrooLWy+lRoS7OkYVF
SDU7Lks0ZSU4QMpoCykWIIkw3jCScm+vmIzh1R9d836yA6WdTGFlaAG6YCsjnGU2gfsohTnh9YcL
1vWL+ezfG08TLqRECoqirY6qvQ3vIzthAEkejI7ThnjKTB06hNsnrl7pEzvdovyVR8a+1Y8Z+TVB
38hT2b1DStvJEvZMHJolhWNJeXs46TfC5wFGlhrUw5ZkWC5d33shsB/NygUB5L7pzeKIhs4qEpGX
l7g2C/AhbSbHrMqUGSjBONKx2EFMedk0uNUjDcc0Bgx85GXlauns+y1CWBXwjB/8JleTtPfGZGRi
t58NWfzWhlLuskjuOTeQ9K3E7bRYmMDVY7QfFVoIEedjQmfYvevdWxR4k0N4cmd2bjZQMXxLqBhA
j5qkoxKKj15q1b/jbhPxlUo5DY8gOke3ox5cOMOwNOrxOp2XMcMIHKJY83VSmZ1GAUgAI1ojB5tO
SBL/x5JxhswrMv1jRhM/R/AeazSeqyzhNhCR/Ly0Y4+FPO8tNtjeXJEPE9KyvfbdKWdc7ZAdhGwX
CIhC55PDbEUAYt017OOeXuvX4RunS+GQTVsKKiseSVeJO5hBOagt/rLCJY2Y3XmdFCVFH3ocR8JA
PunFNy/4J5nPaI9waGFYJ8oThwA/FYwR59wu09QcYboHWfoRQViAIsuvBLky8ujxc1B1CDqUrSAe
zkyFsKTx+IBypc139xnAeBOyFCSGE7xGJ+a/asHDaAo5S25zgipZs5lmq6EmYIutyWOiR3z7YZW6
9vMv09TpP735FDfi5s6v5zxDNCrg8UrpWIeSMZ7D6b1VaqVxrVK9O6616fYK/BnHx8jW1yxNKvnG
mxvaK5hs2CSYy+n3xCDMii9pnpxIkZWnENzrovCqRF+VI6x1mKLYEfmXKlEq5HtjUmII+gw3f8N8
nyCyau+oZJ6zIV4qUE3rDDJbBROzipNYFmOpCd7tQgosXVNTZu5BaUmdWu+si319TfmMKOQ8C5uK
jzNDdWVXRWSaKGnTRjV5fH9e0/gEKMVvryuJkNxC/HUsf3SAnJQQIX9+BS/15PcJwr/owADgxImr
IXiEw277lYppOr5dHrz2uK5mQEppAPAq6KX1O6AuXXWmADvSXcjM03Rlj54Zyfq4HWX87m30qxIK
5QXHy6FhqWq6DBV31vUbt3IayOEeDMk2RNiqFHPMoI1feTYW4Jclg8ItNy/YG/nS+cdcEm1t/RZW
xCmQf82SUBQYfCgD11eoDsTYsvNcHPM57ER3jwUaZdGK8E65YphNnPEonl7l0jw2g5iOggTYjNT/
lu2+PrtotAN0tcDfMR9RyaNFgiAy4IDuOD/dGSY5xkAbaffRBeS87rlufYxG9b3rtqcKsaLeeRl6
nLNLUeSYbs0ONeOzGSLbMNRj4l1gI0wfNOr/I222U+hlrQ3oIyXNjTJout0wjkIbH0NEjRkwGWv7
PeoOnJ4IQsUA5rpkaBcCQsGS0p+GPUCHfyh8TXgNSMlU9CUuH60q+il+TyOrIqaq+ghThkYtVgzO
pvAnaLutJCpiXRXi2Jr853iBo/w3olbOSnBABv0ME0+GbS5oYUco7V5hzpl51ivKTwElnlDLUsoE
LB0bxEabwLUfVNU0VGncRJrfCE7jyjA5AIMIyFrasoiZxI9KTy4vy7eS6vvAe32iFU3KdrXt72Vz
Tm3HIXC1YHWzygXjkg805MRQ8UODX1hxBDukCC0Wh621kbkUbczOYbrpdUXK4FCowKJb3OPvUmIQ
B+Cul4v5aPFIWLe1EqQWXs7FZ52dvf+oZ9zS0rakWMi93YLNYma83Uffi8xOrYVzkbVgqLXXoQkS
a9xzngAUIiajGXiRlBiQ6scBw5reaomFwubkcLXqUJVnJPxce8qdo6FuAHIFkuDHCnR7Rh3tM2Xl
/Uf4+w5fXDwrUdgPLfAYwGylWxRuQXX1vWWjh258u81PCzmVrzKQDqU5Yq4dUKVWutiK8fVzVX4+
nAw/o5vyl1wV75OR/NA45LeXIWS0oZ6gjwG59LauTrISgd8NTp2OnLdYLFCmwhAIJDoPhQVfFB2l
Cc/NanPNWCDV+hkEHK7r/DvekZ0hceYRt+eOl3CjzXJZaG2F4M0KopThWNiAQJDW/fFrwdJonn8i
VhaHKEEK1rmzN3TOCDy1TQBhwDfiQ1UdF+MGccWuP+FJ73gY9QHu2JfPQjJUcWM5sqoaWqXCoxLF
WFxWZKQHP6ubLmXTf35InubXLG/RR/tEkzy7kndtfX/qjGqPHcRWlHT6RzWMmcBJbZW3JkyBVbVW
X0PVb+Q6odw/kmJGqrjRMBgrGIgmHo3je5EmiSM6RVjzoSR+nwZojQnc4IZ6a2/kCBB0ph2BWIa6
lVP4IP90J7qs0kZC3heSVp53wk0a/vvDUkDcuvbHO0PI0FeLc29V7zWdfw79GP0ztPtIg7Lbc+Lp
7gDU9HK76a1Rtcxz7c8Q7GU6lhYin1kjY9yBW++Ye9nD5M7v6bL9WIzJy23cmEObGfx95gHrygW8
/IH6gtesxviGrAtjqaRig9gf7xuPEE5UA5Njd8FakFEIQGuSv2gUY+C9lpczp+QLFK6546PS8jIS
RZxbOWa7KxF1pzvAb4GE9abLUuENi912d7AqMnaQJNL6RiuEgy5+yauHtgW54RXOvx7fQC2aFvud
/ppqwRwdSscYwND+2g6GVBhuV3FwUiZxUKdYNgQRfVS2yKFYktgoQvigJAF+aP42+RAA1968D4pH
qFgdVPzOcv/wx6gPZ3AZCiRPM/nH/JbB6owuT3Or1qMdDJoo15y13R9pEtDIGe0ikQStIUooRtTh
dfVTG18KxNBoq7YLQV7O56UzWyX5FYYCkc6q3fjNoyA0ZNfhKxAuRq2ogdLH3Qh96ra2W+baP9db
sLyAq482ISG1Ir8vsRqskItwDc4MGqEdvWPwJcUZ40DA6zqViTicsYxaHaclibH2naD05jIPMItP
1gy5E3+JMoEm0Mgf1S6yCPCcY87SQRo8x0rpbqUIkuIb1339DYNXRiXT43VJG4eRHbvSSSvNT74w
FmehysTR2+at7sRUndWxJB6buSdEcz72tbkcC4A7hxqkL+06ea2p0DsKroFs7aVg8ltsUj10+lQM
CozNGpMawz+wwQ7q51Buad1lzq8Ew4J2eH2Cbvi+PRNIw96cGMf27fUxVlHs5V12rYb0RQsyn3nK
jsDnLngZU4m14jyjsQrG+4cEPZmXIJgHXBvCdDtCRko4vvDhWa9NjsLqeC30zGiHXnZvKUl+F/vG
73SwNX1H7fd7W58YvK3syev/JGD7Hswn65eLYBmGx+yyNUcUqrah6t3INWGMJqak4Nij2JIRr8lu
L/iuBlBJC0XujzsDyDaTFlWbHf25ykmckQMVWCdE03HZOxJHtFy+0z/jq0SAaquE3R2ZlLCLLiAK
nNOFVdXCncPOCDxpwffVxbmFyDW3ucmc2NI5ciT3MIHeWhuSYrG+vzNgivvJllSF0yeW1gdRd5PS
z8sZMiArEh7Aa5t0jLINUlDFi47u5awUxjVYUzK3oznoG7lY5gjRVpJXA2A1T/YnRSJ7EJHtwo6z
o6lUz7zF4PB1n3iR31ALw4Ooi0MFyv2AdZe0lPDrRpZnJtl+ZXvLFWr1WOQKd6+24IfVu3Fuawhe
rzlzZ9Cf2mQCr3VHeXDjPrr2VTpiaxRXlyhFd/LFk4oSmiNOLds+rh5c0JPpnA/aI8ktwXap1juj
G/DCyJqob1Jp3n6QOTSzXKKQ/0PMcf3Ka8aag2g6FvPjdV+RlT7r/5p/FWjSg0uouQtJgu7o50nF
+8tawwzI2YyA1g63JgxGzxudE/eC7Ag2ey0ymMKFZQacyRXaeiR6qEmrdEFE1e69uWoPO3qL9kSc
QLRB/qXS89tWFfBy/awf1SZEhhyIvIeQWnyNaNiEeIMxwUNwb55kL1ZJRt+9KI4GQXgdyCidmE3K
o81Rkq3jgsIfAt8D+saALZVP5PcH72x4p5ZJc7qXD54TKFqI1RVdb2fvty4/KflMtt5hXBoLWQ+o
KqE30wSN0cnicRntN9xrXSYglYdGwUf9uQNzAyR0mrQZJeiAH+um9XyBFhMiPhkH1nllsiomGIgy
TvQI3Vpx45jOeaL2VAr4Pxcskk0YFcOQtBcd1TtO9jydF4kZQFDY6I5QKEvO9PAOUrxI3BbKRPXw
x1JGEOEF0POmqxKMOHXadb3mklGlQDWh4iFc/K7KOGRS6N1VII0eiMwExOc1SoR8VzMFyAnSCLGf
4rLA9C/yXZf4Z0P2Gya+KHfEMnG0qlM3pHozX1EGA1IaDNiRCvrjvNgoEmryXwVeh7Y0s7ugFTFM
UGfx5vWE8+JBiIUwPQPtxhCytAK6DV0+k17U0XeQxOVRwFFPDfJwotz8UFn23OAHCwpflUElmD+D
pSc3SWZDRiswCYOaurb5mv2RGSPVAQsDrYuYaMcEGlHn//9E6W1gfNp0QWTgfAYHzLhj2QW+UMIX
RZpVgeZRdQjcUQ36nQAzKaAKR81GTfT9J0hJU6ta+R2ysvO3eFqp+fwE0K6LPLARkfa3dF67rbCx
HBWdWUm1MtsXHSVx7T87JGpSVpy/JbXv++UMcuMYhE1J1/Psw0CAJ1E4vsA2PvOb979QAmlvSYSV
XguxU4k89uV+davN8qT79J3ptbt32zXiaM1JOXqNfwjTQwJQdjZDOtjw3z232xfkWLyGPVrAfE+3
kHyrNOGKRi0tGLK+4ymdBL6APxzwad1qpNJ4En18qeHPoeJkJJYzibC7yGsUuBz+fqf1XgW0LIk2
k9sdcAPehOXpWGZf//sGo5Nv5Uq6TOWmnkHkJd9S2bYKuL8izM+AgTG559z8LgPJ9MirBABRNnPW
jrEaA5ixZcT079SL+YmYjEp01N3LIDIeZDByXUiFDpRymqf0XgpCp+NyuIfYhrU/I8m1Fc32hmhi
l3fD/vAJFcA5FgQ9+kh1OaQmlocVf8uCW8hrfrPb7Kz3yKBT6nRf7mPZQOm+UEok5JTb9YRZfNjK
BlL/Zr6QaN0q5B1F0JWgNdhwIFW2pHxRTdJF4L/NlBPbZyCShBcqN8mmhy8PmaAUCmFFrx0QzkSi
LwcSwK3aBmSAHfx2BxMSKnU+wlI/KMBq16888X4otOQUY44VPRXBXc93wFZKrifL+34po5ST/rf0
lcHdTdeXxsltTQDgpy6/G7SxLqtDIz2UQAWoeWCgupQSC6/2q8QUFUuSTF+BlVmEmEEMhvtloRhp
XZR763AhSJeBB67cms8+OMeLavRa5CX1VfG+BalaZY0r8Is9vgQyYcTJbcJUCOIfuhtFdNES6bYX
vQOrGqCo9Q4EEAcarZzoEIaHutsnORzdAkow+ynxX05EApz2x+iJI25WfoK8NufShomeAe00rLcN
+B701rIwHZ/Y07EsNiLxu/gyO7izoIEprH4W1bPyOWMT4iQeZ1IorYbZA97R35DK0wlOVTjOTCAY
hffGj0YUT0+TszmtiOhkXYXtQe1n+SgGVzpo2+iJYOGKTKnNDJ5dTAHkrByTSrjfk9aVWpTThDHl
0ppZQmZkVJI5SpZfsMJYVzeCv90AKAsAyYd6WcX/UTrxOlBwIwJali12L9+FBYpTKXAiAZeFltnL
zMVhN4FsAZXqxa68J5+v5QZCnhYnQTshKjptPhEwozhFdhbfHj5bZuxUV9HQnU7004UxcSqg9l3a
gW4xqLj1nmGD1JEZ9JmaeU3c6ATQe92RO5uHW+GBqU687CtFROeKO0WIiWZftJmFOoydqwVBug6C
DfZcl8uCV9Mpvx2QXpznoKapVeNvQHJeZoq7IZeALXK+6oFtEv9DGQmc9y8sKO1M4MhQoy09QJUw
2ZhrlihQJTQcszZ6PMIjro66IB8ZN+z1ziw4vRGz2SJZkzQ/NxLxTqiTSTIn6xpuKCj6ab8/S3N+
V9l9TXAZKvYmqQo+ralevTAYEhri/7goVXJ2YFGg/KTy0Sse+jroxLpo+8PhtySz8izyL44JNfRV
OoJiRfYEmuu4alV2wmbCmc6OtzAiy7fRBQ4stVJKz2zl3JtoSZb0RZ/ui6FThU3Qw3Ixxov9vGtU
DNC38z1LeQN90tdIIO0sleEkuozK6Fz8H0rhlkkgRt4bHmBOPUTH3Yj2w9maIDBKI+Wmj8Zcnfmv
cnttJXHcN5uJWCMb+yyDUTYnlleoPbaTYbNfcnZZVVCTsnD0jFiHUm9fBpHnuFXSRHm4GtXPcj+V
UlaNljavPpUKX+mrEI0eImmfqLcmnIG+OtyPOzjh0+kpTYEqnbUfcA+72XoK5qUaH+2lYTTPHH4B
ydak/B5iwr1s0B3dFH1sym4f7E5Aa94P7F0u4fiMTj31ZMCxSNRwLJlwU40NDIdaOXyIGQosOysS
SMaHAU0u1KSVUzsacwXv0MC0r572ixCTvvTSJ2dVDx7ZLp8Ae8R6i1SqE3E19OmBrSTva3xHbuKr
f9fdrwy6nLYnpwqR3Sen4mmuf/BIehVAiXPDPB5fO7p1Iy4YBzdoUVz4IQwQVss+PRhzN7QW7ex8
PIQJ2kW/zmqErKI2ZHfb8g+SRya1g7nnzVe8m4oOBsVIdLxeiAKp7t3qeXHJPlsExTwQeZKPgR0v
B0ggYcJ9RRUkdUAo25eUHYHV+8HKTTiNat3x60ksrtbGEDt1HKCrzi+5Dz370XRZpVwU91BEv1IV
zFexy9kpcdcfVc2JUgjg+Kzhe/muasXev52N3T9ZacLQeUQump7yaechWlpUwM26ELDKOUVF95Rc
Z0ouMuTkvUgLW2qOO0d1bjfKdN/fyFZsgKbL2k2ddghOgA6D2wy41qp0xHQbRMhAimrorIboSXmq
ml6JKX99RQmlHByFPYEsLDkjx59T7tpLCdfF4uCjgTWO1K5fhNwUXQqrnBSI5I8HPBaxZte2FwHK
52YD1q+xwj14uHDlfALtLIqG+SMPuJ6CKIko0s6+dOat0cVBGU7R+9l4Gx5wDeui0jbFHm6fEnEa
sPJQyXfKUFfKoOExTxgOA49MAbI7ZvsYSI9JEPKzFG/68oacbow+YUX5AqpZbDo9X16VOf7OxEFr
ZMoNHPbEtiSCY9Gidul2LGImohnkVoJ9JsDfz93wR1d43n4o3Yab9p2JiFsMqgW7QFmoq1hy++hU
Ld/V0/EoFPddNKQtk4g8yrLk1pUzL5rrNPOdNaonWZGBwczpU+czM+hu19WE192eQ2E/rGsKROdp
yiPcs2M32kJnlWWd28/4QWm8G8flrR9vreEJXXEUqjvZVK02QYwezZeNiTqCfhGs237NR/6AQLvE
Rdb3lq2JC32ACYWGg6WDkhtf6C/Ld2GYkzsIHbZyQdU/nuOIbn91orJwue++VLgmbK5cXA0n+yvS
8zR6iOueD2vUr1B2T55M48jt5jLxGUrxPPk8obWCQpXwQQJ678cUQt4eKvSLAJv7NzTvGUMMwb3C
Lzfm7dMuHAHoHTssGjdwbe9lcWipLCZ1n6TMoMps83aEDkyY0jIDz3JHUcdJRVTK1gHSPHT3RjTA
uIP06JSIS+U0qNDo4QD0eiIxbGJ795hDTpQSL4RuC+N/biPjPDIAJwVdQ5KNoCeFYzhZXJsQYoGH
4mSZ+LPGzMDZS88suDi7sk2SslRWjOf7ydPscKF56ReEW7HHPgo11/D1EMz6N/6/wDlXuDogJ9gL
Lu7AzLOdEI6ssPL9mCF3OxF0g3ndxLhmRzZS/fbuCVOCoVbI88DW3vDrht69l/+6pH3eDtLB5322
QcAsWZOJM/AAV7HBVDU+SfOw/+cxcAqzL/NUGP0sMExCb6ExpD5jVQSPG2U62jgGvonSckYH+3L6
nfq74lsTq9EyE68w2kZ4cd9uebcvwAVQ2s3W5sCxvQ1jsv6Yf1nvHzyZJl9k3bSWf6ONg29cLisQ
Cd97G9plvxubPG8wPxV2+TB6WilrvVJ/TbQn6YWJed29TIv6R+a+pMiD2aOrVj/M/tgdWtyRW6QP
X4O18sTfRtEEgtRRalJZFnF+r8BnSp+bDg94veuxFq8xPx/6lbQ/pSEeciMEdvndOf4jlzvVExj+
rB31N5Tzk8JIGI4fKH9KW6ia0BIJNZw0pf8wwj9de/Dba6HfaPu+PLg0bA9qHf/iWHlU1ldGORvD
NhFqV7dw7rAGZUGRCTS69K1lUs+8Ddp0i/23hQTXpr2qWEh2KyFkhV3RydpLEl1yedKyRckm2uka
gECdhovGlmaNp5pUoVnPEpd7fNHjjHcbU67A3L3hKE00YaT6IH55MG+/L43eS3EXy3qD9qTmCfJE
+mASz/5EoXyc0jlBI44Ol4UXr93b3f/gOyMWiCYCuTTMcXeILPh7OrwFeKf5HKyZlgHeCzABZx9W
GJ4f1eqPZproSiZ6RhfIQavOL65BO9flruDTwvu1W2G/h69i0nNB+0qhdZXyQSxJ+hdQFBBb4JKR
PvHpTWC6MWfU1HOE26YRj4zWDH4udXMb2cPYV7BLtLOsch1frCdGF/5UWk4xTtBVQUFgbVyd/lCo
nG3MuRih1Xd8sMm+BXcRlhV4tSyWOfnwvMeH/jXpC1nOheB5M5F4PN1AsiTFx2PdhPKs0RExSi2H
DSghb1kRQHxvhrl1U150Ud/AQ0MYKq6TWFrGpZxPBQU0q4KRj2a1OhjVGkJs7kUnacZGnKNSNeoj
K/tNYr7/DcF2GPVYmpwFpqo4hsubQKt/cnb0K4ljdzJ31PEhclHEAnyrBIDt3UGM5bByM0ihrocm
tI9v2s9ya4hggQIBTUvVwH5QDJeMMWIIXHq991jVXC+HaUOZ9J24u21o35WWQ+pYg2aqlGo8+XZp
v4Ku38FLX26sw2CYRAGTKWEHSp0AXsE/lCOdQiwDSyUL+q9USpT9bM9oDiViGxXZFXlY+uxiKOqI
bm/CAAmd5E1S7K1/czzS2sNUpg34GypWEnheKvqT3jHLk7VUtNnZit7QhYcOtLhpqlt34eL5h9H1
gdaNU6xv7qSDKSSfgKcntRnbLw1gcsWXcV1/dsCBxe3SRZK3LstHfzZtpVUHtvbs87iqEUfFdVdG
e2jbjc+JKWz/cyvkSYfRZUH+xKHjwgfOzUqLrzp9w/C5Y7dSG+Iwt6tMr14zK/hlzHKiJz0i6WLO
A2/DdpuOgA3hjWN0EVzWthlCB8MapA2rx3tSo+jClP6qevc6NzunShHhKa6sn5p2SqanJsjagK8R
Eix0bwrOKBfx7wvy+fN2E8dvyLEiZ1jWkesuKFJL8tHzzBk9s/jCdNxWRxwgn9ucWDI7my1dssiy
NOuEoXeZ5CMaPBgzscR2lAmfbcl4RsH1rHl9nd49qdxmQj6FL0b36advrCwFzSm5B3ticghjWoKz
U0uLE36lVJ292k/igiS+Y0Jz2iVDw3G4C6DAZmsUbDlXMp7nO/62TdE6Qd6NU1KJDSMtnrp2Xd6p
L1Pjhj3FT3NdvPg7tloKDrM6lQZBw1TCdACQYTNqgpVuyRmAcQTyblEpUczwW/7mNgrmsWGIEyOj
spVxDcbDPOEFfPlltekdXAM2btSwrbgSmnVQ7Vw+7PScUNjxq9FauhNCiitpoQNPuYEv44WMV2Yy
GkPUfPzpLx95NpFgBHO+KjPeUdBloWhYnq1rnCRvckH3lfkTHlVNH5TQ/WRTPxzI78VSSZ3rLFyJ
lnwMkIoP/uFnrLgu2ToMCiXR7Q2pD3IfHQeImkDw7qIfEnyoH9HBqw1GZUQNLJyrMqpZFAGWCY5q
mM90qxzd4EfaB0hUEHkWCNE9LewVwnPHrcFfTR2mUquEct4BvsLViEhjPrjItrWnCend2H9S/Fvo
p0Cywhp2Sf+rV9NKovNN25VuxTWwI4X/1OXHeSe7R8InOPU0hmvkVhNeJhU3RmlDikryp/s0XbIy
3xgrFCp6f3KQat3rWWcAHU5Sc3SqOEf8mOMs9PqQnybDzjxNOuxy9BMMxAS9QJXRQtUlOXa4E7+H
YH8hv2hcIHCILiemTm/MH3z5tmXR5G+SA2eo041vJBtrixRFI9lsinjXMPMdbA6FuazAVMd56Rsk
OYqdX6VArEdlBHRlnrOXIJfXKJp4EMkSC9XNVTD+oaPi+Ucsv0g28Ft1lbjHZWv1XEOCcL3BkPZD
R/0RRaQDO8Myv7HKmYIsVwcOpj3os/soRnmEXeAZM7xAatKWZB4URc1cgRt8U/Yyo8J9wUz9L1X/
uEu2b7xOtNFUmEG/NMLDTw5nQmqkKWHIeLTRsrjaROHZawhhJKfk1vaxAX1EGhKavJCz01LzfqGg
8l/bGliO82TClKlWshXVuBgjl8Q4ig/ABzrJOBYcwmXiArdj8NC8pYo2VPU97fjPKljq79tF17f9
tYoDY8W7x67r4uv8iRyNi9+LdvY1hDdAIc3rg0jxA7b+5yR4Y9RTgVzsyBAC9gdhhymoPEy2CcUx
m8t7mNYMVsi4k7s8/ejJx9jgnM1MJFOQ65dQ1Kl559SQHD8GVgALl7pTpI2mCAlh3EJyjK+yS6IQ
kwxAAy0oZrqGs1FIO63CKQ8bsTfFoAOgP8PrcbEsuqloG5mOc4kGfNlmfE3wo/l1OYdfGGLeHlgo
KgOS1jVPdzmxNVjaU4jLkIhcmWty940rGLoFbZCvu+ubWKMjz7IpANr2iJ6TtufPHcZckedT0k6d
ykyK3M1BrxVlVeWH8At6n6ovxN9YtylIjtmp7YNH9/jUtCRKbL32GRchX088rbsc/gs91n79jyiP
k32xVH4+Mj+zIiSbozJu8nJ5L3rVjA+C3QNGjPYbgOwLL5W1RtJZmsE0XbWH0VtIQbYAZCDpc44e
cylissAFrBly+OsA/Ck4sx7b/Ry5WL5vEp/ryGn/BY4GQN2vWrhzSDi07sYAMNGy7AS7p1toZW/h
r0LBmfaxPxGVIfZNFwtohAI69pCxZeHKXMlxprIQWS/4zqZyqqXaArpWlNLLwOClaLzdLuIXzy/s
6TSZ42Bm9URb6rtxYBAfGczv2R/AwcMBsIh6CMHIb5I6VRSDcgSQdDxjRq1LtcB1lPbmobnoxy3S
CCxAZgB7n1qZDnXL+aXPs/bwWlp6XGz8NsoP23RN5Ad5BOpM9gKCZ29dpVgovlONLcV/jB/wr2v+
LEI59Da5OX8yO4mcjusSnNW7IZ/kt8UNWt8x9wEkpEymcPcMYAnswFduJmLqCUzL1uMFHu/hHNB6
E0AuUXVJgOj9CrQwDqidRXgNSReAIYzvnDIlUWHcb/XcjNult/Wa29+n9Dl/v0N9NqSu/MnzfyQZ
WS9uWAqSPGjdgrSUraGGODZwWGzcxshy3Wos+puZBDHymH/x8UxQiqlTlAPZ4jNSPzK6oB1A6E6f
7TdAySmYtwb0FTR2mN/p4JDinaqeeC9tDRxmgfvBBtltEgPta/Gig55SxjpiGCYPjc9cqiyw1+hv
3r9er9plw7txJY3Updje3p9L4RbWiFOKkjrkQD4TKRkn1397huI8Sr2wZKj1JkC3s3yqeTfDGGbc
Y+UFVmsHGR8U0IR06kV4J1Rk2nmR4406De7WUbCjtwh5uHIIZt9GE9yz9RgaOM65N0uOyIf5Gm5l
+0TDVNhBx+8ws0qCBq231w8i+EMSV7wV69cTSktKGCyFanFZgRdR2I4gWuwgRNtHO6QVpSIm0Um9
EobmkAL0siQ05AAf1/bKrq+cQifQEPl88MHgbWldjmOKnogas5kXyFGrLyfGYhN01+WgHMPSRHki
lL2D/m3inTyMauiOQrfhMI1BKEH7zUJ+UwIEuLxQJu/FbBTfSTwoANfLySIewsHnlj8b/xvJuMZW
4niwfju1Tv6a56lCaouMRAlBwqxdcRl1DRddVWL2gAM09ujuWnrGFB1G7sM60hZ6ObDAJ2q+uxcw
zryFPbzY5aGp+WYecqLGt6TYlMILns54LEfi7osbr2Lgv6Fy+xN+/WyeYt2yNnDvzxyDt5likYXQ
EpGqtKXSM5TTdbMBzGFgWCYJ8IOh4k/83spn6ik9pmk0U83+UdWqMm4dcVrxXZ6IMloBJPC0lJyR
QcXGkbAd/ijBkdYdAxZl1xH9yNgFUc7/zELEWvfIHwxPjBQT5ER0RWiNeeYfYfFshJDUzt/DOCds
E49+dKrxVsf7tGclVe2dd6GJpzJDQuyc5pNOT0tgdC2h/PjUetyZ0w3AnKed0oYPIbqItRSuPw5R
ryNzpUQPnkyu2Y9FS+2D2f8Uy4GARgrwpqpAOD3Skk1FEBSqc3EyzSML6eRucVuUhjEXzjQDpcov
Z8+zDUNy2Tnot/k3Ndx72W7Ty6I8xF9Im5ZwGDXCL9yhnhnYpVgL6hUFlAWiMUpF4hz8ALHehQn7
yFAzWg9GcdcUfIVPNK+454eNUQYFoLOFREJ89SHJ1mx8PRXBDZcY2A6vqReO9bHRwyE0cJMD1B13
YZTJRz86NccD7yMyyTi1mHmdboDIizz5G9awdY+jkANUdaJyAteHnctMvQeUYcEg1uUd9lNvs4IM
aU9rWNMz0UygRSsqCp11r56nGgQwjt2TqiB+F+p/R8ARZhbzcNmPWHpJOmcLejPB418ADWaTBnKS
2RDUUvyIDixJCJIkEO8vOCBLZSEld8r3PNkXx3qn5ajhhDUtHV34F8FTklHV6x6Vn+0JTDf8hcOb
5MiWSrAVUxZ7mk/0D3qzbNjmGEQlxyh7I1mjmR0BFzy/yG89hvkfQ/zBk0H93FwYjrFVU+rUyxeB
MNBwtxIChDmU9ltnuu5RV5DHC7qC8fwBfhpmXgakPqwaKAD7aFQ5Tbv7QvfmeFdAJrMhN2cnwp23
lS2ddDPsN1A4vNEcWSnBemXHHJua2BLO6IaF6Q6oO//sESpX8ML4bW71YN2VZBqivX4HhFEF6pOt
nGXLImvBYxh35uREBSSp2EbTtPQMiVHUKYPAEKbRnOsFLyTNAWZVYQG7yIc8UFqEoirpnO+789eG
+Sb0bm+WFjSEBOa9E/cS+vhAVVnItlqqKxyUmc90oQt9OYEUf+aZsCtcSzVAdw2rpRmAEK8FVDkf
cCzx4sFzQqNT9r6MUZf+XZuBFhKfZEaaWtVXgCuY/nI9ansXrYtElGdNemb21JF5FRJZUt1PEHYk
UJPzP8g1M0wYxKhD3HEZfiprHhg2/8qoFCLlHpZlAuebFwYi+tdhUXXG7mGc8m7qHgwb/Bk/ZDgT
nXMsoRebhfLZWaty/W3zoEjiuoQkHqZ/wCpdHWDQix3aCg+ASoJ2fkQ0d5odzQjhUcwzXo2fQfgF
NBPJUrwWgIQ9m6UIg8lFAfrSKgSf7oSq1j2OgcXi2XlzhB4ve4Ki/7cSvIg4fP6ZTNzLdnFbnOzj
mRnhmp6jFCbE1Q0IDIw/qySc0ZG768J9GsOUvizOd7I22qrruPk9NYtBid6bFSRa1Mvf5JN8GVv9
r19kZUhws9kc3zj4/CkQUgWIt91ubu1XZAi73k2/fT9b4LzQS5UWsXf8rccMLWzMa1bQf+H+unI8
sCbb/qtxReAcLvbwI+OyZ7wHszYoKcVqFqmL92zPdanGfDM7U5zGNpWXb1p0bcUZG2Tj+nDMNf0E
0GKayvWSqEyQuGELWeuO/UgrHuX0bm+d9fQqu0c/5UbuEnm8F3JWgpcSng3yjIaTi4lUR+S0wQJc
h7rBV7U7cbAcXurMuoGUhxxEStRlJ0ZhXBasY0p4uI+H07MfM5VOX6ppWver+jI82bILEGglEsT4
0ggc5FDJJW1uG2UjYqlhASB6Cn//bexMGqn4jF1B8L6w3szrC2R58Kw5J4J6dSbhvCc4ZrUuLV4O
9LRO0gJL3pZRJ2DwYnxGpttReRJGvqEmL/rKvPfQcI5bqK44KsgWYdblZH+BNyk7tyWHzNoK0KVS
lMq1Fq/OIrblbBpfLO6QBvGGCGk9NwqW/nowblWU7gibioCtB1AlW6FwK0EcEHwzp6YqQnUIikKs
5ccN40BeV7THtmaWkXGacZBiAqaFIXt9hHdlZ0ZBXXxhhnlYVqwIso5Vae9Lvst6ufO0RxHvQ3t/
yrBVHstnv5wZFm+fvyan6BF/8znB8k+gqTC8ODtEsLLLML+TbGKdRaRg0kAUVEXE0deA4SUwZIw5
NnCl/tgCUtNb89jrZpP9KrAeEJBKB2aMdgV2QE9YIMudrL7xKc3HmihUpRxPjQ8S4XYiN5A2dVUD
yOIWEWoOTI7RLlKNAf5dJ723sVa3VIc52HjIJRkV/DxMuyij6FjaKl8UMYTGGzoIC3p++k1harVz
XP6CNqrLDQiGJ4gDpbDV2G7V41SWudfbRNhhJSGpOekuL1PaIQ7tj7CkyXZ3PUNuhMJwXFHPf4nf
YjdBFKpupmozGjZ8jLcSJQViqDH2+G0dEbkhntG7VDVOe5AJmt572jgDaQpTYNAyuMhRYFdxxqM0
HGP/1RTfqB1fLdOh2i1tvNBHT7mxZzI1eiAp+6sbxaBV6sQLQlMH6UgIFzlfCbHLPVroi04bBODA
avwHtg2voQfZPcW46E8gunuHHb4WhjeYXAeP5/UT5yTJ42d/66Sq8zsQDDMK+hSrF+AA69uo+Lc2
/2IEp4zvVW9oTQuuyFg2VHt0gBm/GayK3tjhBCbHsIZb/+81YxGGc2gesfUcfmzyA4dToy+oq8xu
VTLaLjAy6TIMKyhm6san0YXh4GO2RbIKekATxgx8IkPQBCaVmarwHwKiHnu5ezTUHfSYUrik1PVM
4E/dldWCh+fr1hNfapxmfkuJ2eXNvUKwDW4JAtdEzCjAsFVUwxTNy1k2Mm19fj88BMpFkEONuUWs
s3qG+43/L7f1yTOFT/GfwAy8krKuRD29CKaTDgzKHp+wNt+/SHAk2124so/fapmbgXKV6c82UkKE
6fsA+6RdmCZYX0ObZl23Nol2cXs5q6Bbx8xOEq0AU4vi0K+wMJBoJW3TTs6m/IlABNkT2aVJ6Ufk
TUnx0/bvvxc6VY59O5c22453zDzvTws93m5F0HWcKDuSUaj5LqMyj41mc3hNOEZ5lpilM1NqIoi1
o0NHRlr4WzudaKqqifFNU+GKV9rartjP22n/HEflHU13Oa3PHTCWwOPFz8biMTM5sy0Bx9kEigft
GAd5aaeFIfF5QMUAogPgI2IGbARMl45yYRk4D4tteBHxDVhRIArs3A2GisRV5s83v606sDmSVryd
BTFG2eJSKcAMrzRZfsQz7XDPuOxK/BTztVqeXIzIXQx4p3CjPQqMaNYeVfU5BPfprjEx0v0aRZD/
n/NaslR8g7layQxaO6+o/dsftZlfwXhVgWtrHcIQXI/4hkbgUbQ9QVtSd39zyFbI+qccHtw8EOu7
CouwX6dhEElQCRVpLNb78q4N/iZWo3sohZ7czoLmsRpG3swIqxD3RDPnqm0CzsPWYQOsw+IfrH2g
Yz5NSMwv3Ju+1f3p9P5uYycWByH/K10rPR/KDltP4z8kZfw5HfuGYv70Hjg7VBTl2F1tTZUjVGn2
C+0asH3YBGy0FdgupZNaBDCEUsK2a9eHNR1tKTY7NojkbvP0/XItSDSTZ/xOnKuHXk7+CrlxH+jf
xvQSkDOTI62lcNUHJifnh5ubHxd7zySjZx/Sc7eawlJSlu5pM8Vs9ivN6Rj3B21b96Y8TaANq+wQ
kRIWtuKu1PEspNy+Xxouraid4TognvQFcvKWAOF87zDj7E929vWDONhP4tI/SU51ew+HowS1x/oF
FefX75K0MJHZEMJHL6hqAUYbBcxwhxuUqnId6nRUWeQ9dzLtXuEcCiOXfpg8I4+K8lrTgCd7xZcr
cZHYjp/CbH9YEn+hxcBxCSvfGXx4Bh8qzI3muziy6N/XXIXYo5uSdDW6hrZ1ti9jLJjm0oM8W5JL
wkl5fJPfFJHnsOyU+uVNsO8VMvVe7yTyKIJVYC0pOZ7LZi9eUBrYahIt+MZ/Hdx/DqLjXUb4KP0G
21OmRgbaMTlJt0BXM1T9jn4tOFhZaFtpdGVlC+zU0V0lueX/nr1VRtDRzuVAZnDDGQpYUOWZFx4/
/DeDKlAOLd7L9+7qoAjyRcGs17p282pEWrJO7Tb8xlYvLwA+87kqMTyXUv5DyfxiDd5UjnS9SvWD
JnYMgFiDK+gsbRXjTn7MFOc/1OvOvSoRbyUm2/Ff4haeorjq/d2gGs7qlDeYl2pQUqazhOicSyFq
jhvZ8DbeqGtsj1d3OwVajzt/NC0OOSVYWUStQlSMBvevJ0GHqBl6Dwskpp2tDo+dc/vbNQL0WziL
gm1e3Nbgk9U2rfP+ZbcvS+xfpaDAPusJogLK0gbxM0PU3oe2cHb2Uc6qFVDn2Qz9DKW/7sJshfp4
7K+HCkQc5Zs98qsinkN6VQ/NtSWG2wJyRliSDYPfFJeNc8uM4qPbhcWNV+TExNadzGc0eodfTo0L
J47T1KmoscFTW7ruUGoUaT5papYy3aNW6ZPOPvm6uxROn9rizOqBIIgDegdiIiey++08Whsm+pL1
NGsMVmASNtjrThKZFm1wtu+lm0tBjwlwF+Ktltf9RYr7vBlEluM61BeQEgz4MgAeeYvMfj3jjkqB
6IdSJr28Jmfrh25y/nVDZf5OPGpxyC+BvhJVqCYdcwTNa+ru+87XgIfMv1Pl5jUnGaZpqRa29ILz
P/gsDJaMfTXNfVNEH0agcwxBOcsnnctMex6h0sqTs7X/neKVxwhqXltlFU4WlPd18gbucpMCCVhX
GxGGqNOj6dKJCsv2Q8+PKZqF7ZpebRDF/v21UKYMHziDnOnCkMcYCB+K5SRDlG1LlIEsLZn/SGIS
nzmr1Ja+z/kmZp/W/ahnDbyaN/ZsrBPzbvUyn+ojwsfS3XS7wkl23XdBw730wNJnmcwh92f8GeSF
TYIt+3bIcxATwcsCZplKhhmhKsJUeC8sNLwSoAEqRUR5u3711KmUvSPKiduIlhXkEL5nZgycqWYC
29PNq/8ECtZN5bOtJHTv5ouVUxTD4mmUZVRRRx28DAhCj9FAC6PuaPxdaucPrqt/rkwQkE0r4n2l
klzdrVnvn1RGF1JrWMO+77nbzVgk80DWKuZWCTofD7N4+NSZspPXwilYzj9NZxqaQ5FeyW3HOPD8
Yu5KPFpEDVFmi3O493oeqZLyMjK//3iMpt6moBpM9eHjP33vnKSsFTCmwhT1uHjiE1pDivuNID8M
FVwQITmF2z0xW7xCnnDdlfVTao6hpnEYldqvM8SUqofECy0Q9D0DrLRy/aDDwloZReuavqbr84Zk
skF1n1CW6fA1S7bYgd8nGVHxMIT/UJ4boElYMapDFE1sFr4lfLuOrllR//M6DGb6h0yw7Yu/bVyZ
4Iwua0HZCJmZUVYg8UnUgxP5tRSCy3VryfzzUvUJBIFSgVJMdWROo5bWQeOygcUypJOpCG/+EQo8
pc5H87H7xSfnQ3xE4rh3jOFSHStFWgcSgE5Lzkcgq56+CtVH6foZGm32Bf4IB6UQwVRoqXZ2v9/b
HtcyQfly1KBDOlhx2s0LecO9aq33O1FDuv4U2cDks9Evv/nWMMVOmrhJIVf6Jkm96PKQpJeBtLAO
JQohdeKynrnn++rpaxjA6XziOnUc7/9VmPbVCX351UagonxHkPivawHcRsGrmf8EXkV1a4IO4R4x
SVovX1BkmGDwGjtiid0uAbK4kGqo+x3jp093tToyVwbsoNOj0sRUDl8lIoWlCSNHEoV5ocq3zmGz
Diog/3xWlV96zzhaQKvZSCu/WJYTI0Sl0HZvhDn5xOiwMerZSx5snDt6gYzSnnIdvLNynjYbUVCW
NHiFv0yI3yySpkV0X0wua/4lbEuKVNBxrtmV/D5HmUi3c8HlXJ139N2j9NLD6jotkzqqpMAyfaDA
z174Bb2QJEa9NQPCKJXwRELq1Bc9LkYejfehPpa/4IgEiwpXdNze1YiKsEpL0SprSrw1EbKaJfp6
1/BGP1KueQR8OhMaq3VkHEVjsYpaK8MSKiqPrgmd1FVnrRJy+w805CUWdFg4mcn6chE27y09/VTZ
pU10gTRb2qnnC4RYxE2Khb4kpxlUJBR14SL63tlkZonpsQXUDLtKKuI8pO8sWjR7SVN3kG9y7AJv
afLgw/jOpDNHNbU5YV0Ewc+cSyC/xrPedTIJyQiXS5KxeMOiA389hHGC3s6run4041WhMlKrYMrG
VO9I68a9l/W7e7dGGkHXuL9rEbVm1qXaPAO1zS/6omEeJY44y1baMnWz/plarnNGn1x6vu0k9BSo
OQ6KQ6IBLIG6EFrCvnWRXT2A4LdiKHSF8o4UqMcLIwjbZnW9dZ4er9YZWdZN5NkAWbvxbxdIiyKQ
8pq4e/5NGN8NTKmxCNLIkX+/c221uekJpyyCHwLfLrTg19lSIBVwEsJTAYFT9jjRt+2dqiLuaBPK
NOni+i+iWQ9kazClkFjAInYWAVsZYlddWkBcUAh680xkuD6hOpoxaGM/PvfUqyONwZKLRranVeyn
AV7XODKRgmaHk+ug/RktTn/zgBUG9V+e6OxKnPz8l+ue+jK87hUssgyy3mJ+WYsayUnZyDP+lMhE
wsoPjrq0yJzQg6B3WlHvvahkUdpiB27RCma0r6e6q2Rh0xbTlcW5dpkTyTIoqanH23LFUvdreo5N
bDv33lOfERtH4Y/05ETFTCXvhrMLxqgePjlil0xcQQSKj3ZlnDi0rxvOa16oC5QN3sEsTWpPrVfZ
/q/updMruDQkxCN9AqTPRNVnSkv/jiTXi0RaTNohSwR27QwGvC/RT6ymKKnr7FCBo0xSWhLalpYR
HuWuJEKDEm6Lw6ZdzoBrBVkWANYOAznF+UpXfVd2hIQ2AkW+Mr5GLXscpi+wcUuj3vEiju9I7xKX
zTcu01WQecCvo/srCbVB0vGgS5pacArhixlFv/o1ROoEMdDQQORgTp7uTQ0Xn1jM/+AE9oCu1xpJ
cTygoqC6znCqkrGPrSMmTihlclI531IMkOKWnWTctAL2gusiFtSVKkYJPf8a2RZXLKVDdn4P5fPW
xk0pP/ItCLgdu2+i0FwD9bheSLOtwk7g4FkLVAztiH9r6krxOPHcIHKtalmu3Ki/z7yshkiQ0io7
iaLaf1qnzy3BFG6LMfs6CLkCGZ+zBJDs+YqSdBqgokE1gObJffTAKwYdcsUtng6Go71c1sFJs1eE
ZNKEIs9VpxTbEJI8zE3y8inbg/RUG91K7WFumHurjD7ADdgFcEmSOua1/+vsMaOY13WkIKOn/LwR
VkFrcRj9loh5JBi+yUMaix7WLzjS7MxOH0VSySIHrK9sYzkaMiBaJL4zBMXjarsbFsury9Pv5kDX
AjlPfFfRcRaRizzEZrpMLxHVPuMrU40v23lV+wQTuOK/ZkCoJCIvt6zxx09FXQszDj17JgS+TzpO
iX4z4a0NG3b08xE9i3Cs4XIAhzRUBOJv/utYcrp9jcKw1m042ehSX3ueTsz/p/BqYNMRoEEjFEJa
nZtpimVctz5xpwZWOrG5wAUuCVyfhb1tHpH6KVU6V/wYfHxnYbljmAu0SBTyxzoLT2Rn9watSlVz
bMXPuXdALPgK88Uai9gzfCCz9xD3j0+f6G/jRGr4K846UZhba/+BwWLtdL6hwQQAOzppQ/8ngVwe
P+r4IFbgdQ5ze952ER1DkOL36stM507rk6SkUvjZicb2Zx7AsihNoI7CTatJOXyF02QSQgtBbXqh
7VcR+D1+OgGASIaa0K/N+w5MylSNGIKkG7qOJiNzAtcemW9op7ec8YSMjWph+5brLBOH5yFznAt2
k/cV4ExRNRpQYMKnBv+EUiqDdOICn+56zE9zA/8bGIciK0eck90SRB6qBzEAiwQ4/poMDMeB0lbh
hirZpXUftkXnDQOrcLVbr/sJI26VY2a+ygqggHTc6+uYyOKaBBb0pfoHQnvBZ9MQEAx1glrn5zXB
zQxths+9lXa/JZniqGNrhl+3mmhCfLMHh0lu7MNL/0RRai8MOXZh6b5JPvOf+4GOwxcunhFT+IDb
fdwUG9r4wkzcXZ5sKeunDI5GiS+WEyFco6AfmiLpg+ekU8O0tjxv2nteZu+wd81SbXEI4zEkgba0
tykZUoiQfo/mDW7jOZ3VVQi7wU0BiAbYBRlJkHE5llkOvMJLoHTmVpggoLKWTKPOZlG+xCrN/JK8
mVR9e/Mb2aoSzaBV4eJy6y+VOYYnXkOoD0BryKVa8ifQX1bBkxqOUe3Rb29g3VmXsgq0Bcbl0Se+
ks6eHm6tCRGpswMpcF4KTmFSGTjt5DpBAYhb3nH63Iwrsfa17VrLeC0kzWmtg8EQclvC5E1AnAAu
AKV5zqTvm5HuS6SEDbSHmaTvY6NE71YVmlZx5Q7pBGueGwF1sidqsVBN3P+IA4ncPOFDitRIiSwL
xhgU00XYODkM5mnQichoJhlOA9JPj+O/Z9OItxrTozaWC6H4kue858M+LJl/Pqi81nmMW5HEd3c7
R60fj5KB3ywiONiYL2tOPIpWs0vdX/NS1dxPOJ7r6MSP92EA3XBaN8pkA8CGckpHX/ZSozzwOSPA
EFXRohLTSd4nyw2aqCx4OhEQLUVSoK+dFpge6MozJiQKttW+k5fD6mQS1Pk/OXDdzbYZReit11w5
ztmHgZCOj6wY1AZZE8jRhHMNxE27KY32ZIsy93t0P203qSvXQeNNvvdSbtbPl7F2BV++MfxYXzAX
TJW46D1n6lD7I6DUfnur4V/NRwwuuNTX8q3xu7uNAXCecbZZrgXxOn0gN8ZF6yB3FpV6PUNRJidk
OZCJcyWDzxjD+H+lyarifKKeLqkUbLcixLct/M+cfcAHTO6THSh0UAPNWRgrfSoRyqCCVX67maDB
NVjhGxCYvtTIFq9fJs67yHxVXU3HTDJBhOLVZfBAJ8B2BbypFhJxPsQK+DuyweKvUZa2cOXDEqpt
eqAiVID0mOiYgkNfvVNRHHtawlfeoQ5gIsd4IaiDNi25AOpiPuk8Gp9zupQUDNGBXsv0YK3cyV+6
NtTiGVRWGUZDaXrmLMFAIpr634AB6beRBRrrj+LrMBC4SN2ouT+gjMiERfdc9xNbNlx7mvnhOK0i
6MYJM4VjlhIdgdY7cPUEhD9xq1hqDBm+hWUn43femSYmaWkGaRIQTPoC4Lz+bqjYpl2WAfzeZbnO
7B+a+tidXfHDUmQbNKdqozCzMyo2RDJFPf8O3hWd4YfOyYtzQzG7qwyB7HBjAGHOeNY4B3q9597A
n3KWLmWirUPSoRCSgvuK71EnRQZh2QITpq+81WwyDnB9UVoNRpQSyt2OicBU1++uqu3qUwnhK42b
GQlwPHJLJ4Cg0iGN4dZNDQxyNAlWuv+SCEoU+KZ2bS6be4ehX8/AXqLIm2Ci46YuwwhXV0zGVRPN
wUc0HukARvuWpdqLrKL53R+c4umfWjpLuEC150lELZuZXiukgPD4m04mM/U4+fGVszLJ8wOVD/8k
vAHQEGV2Meg199oIR9MvDcThHN8oUBEyMd1v8tXw1laHfibp0LK6YOFe0OVpgz3A7WrFXMf5ap2z
kSKphMhnETnAJJGvY+IY98sQQMQ7a11oGPiSDkM1LAXbIFQPIsuDp5BmTk0qnQG4LfO/t+wwd+HE
eji5nDIzs88GI7lMae++/lC3mZ7IpyNn5r5jsdUxen0EkYkxSO4k+v0c3Pm40RQF0NBhBp99YyN6
zPrP7G7JOdgwjg93+GrNNikD2WHCYH9iCKpVgZbhu63wg2573y87GFKzM3/g4T5qkYrePxULIwtw
907M7SBKiMW2qafPaSvigZNRzOlMV8r9fFb723gW3tSdjuyBNZhaLcD5grodo0rnL2Rl9e6na2g0
upMJ++qLUG6UMQ3X9aAlbXuxCmL+R2c3292sta9UEJQ2vDQAEEjiZlPMNFk9tfFk56G8xQvBzYWM
CgRPduGKiMkJxCxIs3hlrHDDGpajeEHEgJgM+Xp2Gkcw+O7gN4IFXAPtwKMnV6bnF2pvMditKZcz
ASp33SYIGHgjx4nv+I5SmVS4foJcvfsgAC4kQLzfyYwycUMox3wobBAIp57KQA4CWT9Hts9xXDcX
qHtTLveZH1ap2ud+96lpOrRUqqRECG06ylOPs5lgZrxXa/ySSAjpd5LNj7+S2WldbZrhcLl7alUR
FjFwdNfkSxnWMjvx9teDwNpJVVC7XJO2xgGgQl8ImbTgs3HlWTmhJwiCAdpU3WJlbr04MO1cGDro
Ghlta9Uy5hn0IcMgtm7Bsc9QVF0ro1rlgKzLtjypqwFEXiHMVopDpYNzhyO9A79goK4PDkqnMjot
NMwVgq12plJoWqI+7HmWrkE5U8wjxBmw12d4XILUDXNuc6UauOz7bw2/rUd93WTOG/Dcr8kYGkEJ
2h6JxoljhViPnw8dqxmLE1Ee/oClUfIntlItic0h4PDpc58Wl8VfcHuHiaupNJCcxHIzI9di7NTh
Hq2JaF9YKn4ZjK3fXr95aP63/hHZdLW/eq1p9s10EfR6KqGkYcsKMluYPsJZi+IDi1M+xyjwix99
8vwv4rFy+Z39ROv5tltJCGn9nJlIjZ+ZsE3+GHutfc6qwS3jqwamTZkhFC3cisKGSikR6QDAOg3R
Gr9okVhT8JpZq0ChutQfaEXgY+EtMx1JP9JTqBPOvXbzW+w+6OrH5hIrViaEE22ljRPPKtPk6UW7
kUkkmw13AHYzADYKenJge13zMEF8lCAmXqB4p1UMu8zOAwxsyBZDkqQigcw5jqi3Ldt3jWWvKeIJ
B9Xk10N6K59KIMhGJi+dasDd6r2Mxsc6zd2GlVuudNiUkYO8rmTRHvexu3JBrkjrkvG7lGANCaZk
UYmuHHTHdaTyO1ou8pc7LlPJzL/ChRZvShMX5zAE5tqTkeOIU78PIKBJyzOQwY9J8QF5dQ+7Qp+h
3degIu74+pFq5V/9FRSL51YBg/l5WJNuHLU+W5SufkH9B+dRX+g2ctju/dbckvvdMNtqr47EQrio
DPY98NlT3VLjDNL0u2a3yLFCFWtjYvRgy9PJTye/C88iNT6MN4FC1pCxCphHceQpEblosCJH6EuC
2I0r6ml5Vqo3hVWyeLT9Icf6nwmrT/c1o3vFf6DC3hZJTycgSECF9No678QLEfx++2qCtjWImYhx
Oq5ZU35aKoKbN8ttyIVgbtvVcCrpa7nQ0rC13VZ8RY9bNY2BEmONHtLYkgJSYdnI3AJv4pSSjUMr
vI5EzS7lKBO4ZColaBFGsRHdTwe8BgOYPgA2gyChkUxyk2Fe1gTL3Whgp6SR3qv2XnI1lL7RBlM+
Vz36P8pkE+bSxNDl0XwngORSSkHm3sp2fzs+0dN+A1OiOUvXBZRP9pEbcP8G2VqTLtL4iQ6h5t/H
KSyiq4/bPL8L80+FVKf5V2gdaOcaYxf03zEZE3ZrIRj78tbmARsru4ZcpzEPE9+DmMezGkc4UPET
XhwoDSmyjOMiobKtgge86+gkxtNEWNorMQNWqXN7NpDPFdMJ6cfyBWT/XZOaopqTnpkcW4w+VeG9
aWBvD2sjYFjAAjH2Rhr7F7msc2Gklrp96lw9s2JNyWOdlc6g1Z/Q6X/C4TYAEBgwzX60OAJx9N4b
4P8NIq//4TPaLBqlF9+6s/NG+xfroc+WTW/s+fi/LJKpJ59ns0ZeVDrvKV24EsRBNlTepWBIAhpB
mh5hspffpHLMEY+GQOWuiHEBAt1fyMKA7nQm4Che1bzkR+VA+/YxFqJh/HJJlVKi0M+NJJwcAWmj
ihB4g7Eefc9cVfSvuki8NXHVF9zSqoTM6I88hWCHeq+nTEIVhI7GPkApl4tLxONSiDhqtYjO/XbP
qpPQW7uKkENVEF1A2LeD+G3gUfizyXhjKzPFAWQZquuSSBn+4/uMVTiu/9VSoNcrvLjLhRjfTH2K
99babhqsGKJn4PvsaBCGm7zA08NtnorPAiHR5izC3qabI1f47zfuytvYCoCyp+aPAvsZkCSD+OVw
VEwidEIHeCuSNJ9R4WnABGztGmKIBCt+uslIPJpvcknKlVWzZF5PVyiQl0Hr6sIeCbVD54lu+u2W
48SMjYN2F7mtEpw4p3iaFCdOu3LzrGsucJI27jKXCpR1MMLGxoorUiJuMsMh9R4Fxt72sHlv523z
/UEsf3Omvt6pJHfBADQf+0yQACnrE+Qs7ZDFUZnatq0gpORc+RADdt2iSkrApgJhgVo4hs6V2j2L
GBkFgNzVlwII+TPCF3q+qJJM4iLfC0VPqt2O6iQK65agjEIphM9eByddcXTkMGSS5WW6/BHiLjO8
x2TIar6XerCZsHSPQrMjobSF1r0krDoRXB8TqjjEJYf23D7QWlEwV1fUEcSnCQ3nPWagO3YxQQz2
Qw9T8eNov+cul7UoJf/F83/VmnfLsdZO9ZAYDw8hwJeJWrOelnVwOYm75hkzUP3lRU9KXIcQYxHA
GDv3ndIFHSvDYpE/zPTPjsu2xM/ZIQg5wtfbGR4peDGQhb/2ZGPBS2rXWWkKnN80jJv0M1nXkdT7
8ECVggFt0AWjSBIn0Bz7gCvBPwO0OgI3yk/s4y0KF36iNEeEHtKt7gMoiAxB0tuxkXvYzy32umbB
FEi83ekaaAtLAI6YIGoSyvN5glOkzHw1gEJ8ajYDvxROQTOtYmJl9Nj8ngzIKEVQ/BANVmMhor12
0CaWLje+ZA6lXjLXGwR+Xn+R6qD+pTa0+Hym9LlWUBof+NLLdqqNFtbTPAKpfGKf/oCik36NVlpN
Gn3p1xeJ8+e8OH82unYIknb3jmH4oaqqYKudh9A6XNr16lQ3KDufIHm3FHIsfDTw7Bj/U2luYcr5
oBbLWCsydFJcjSLDrt1uDzXIrB4bE8p/8Jz93gceWVpQPX4cxqzTeSaoClJZaB88afiOKOWKb2yW
+PmjUJJo5Zv7bp1v2mo6GjbAg/QZB2DZ/iqrk5AAwW/FFT3QDvb8VL3jOJxxmPNLBpcAcYQzjI4c
trfhNTRytyzLL98yN3yxv4mWc9i4AzGNrRL6FfybIp5/ciNNTQiLc1X0bYZbVPvES5lt2bvAjdS2
sDOxaQNbdBz/U5Oy1H42sdeSBJuCbvXB6VcNjp3F+WLpX8x+l3t3xiLvvFy3b1k0BWJGc2M5DrkH
2dnfVPWZIhmfN3T+BvBJzzRJNbWaiE3nApX3aagVHVk0zP2Sb4sRWlqNicvBZ5ejYj4PZY8HkTCP
IZBUq9Tne28gw0StbeoMnFUsjbCdILWRvclaiZ8GjdAyXAGbZG7BFbDjJqdGYhG3YZ/fkjlrOGMt
h8aVzEYY8G91XSIjAeQ95lm/jsu0faiGtesciayX/9xuj40n3sGv6jtrjp+F1OfZP8xmkfTiN/Ax
k5fNKHDbTTMzVVk5EUjyqPTOiLuu6iMsuR9z6yp+i0jU4l3PPlexqts1qOrC1Iqo8tNXut77qm5e
QudJZ9VAL9/X4lcCJY+XcmY5wP1U7qU+JsreP5zzT+9nUcCZODJC8m9qtvKRxO/rkslJwkw5Yd3Y
29fXwgEaDXQx01TXmcJNPqgHNOdRhnpfFp4bL1NMi8J9eysTfjhOdCMwgkyEPBkJx4Kw52twvZvG
GKJUlkwQCIN7/8xZx+xjYAUg9SoeNJSl1i1HiPrPnSbXmXKxrnqfOyRLp91zWPzGIGAWissz2gHn
kjR96i/pH+eSu4WST5LxoekUHmHGRkvWdE6Y7n4P/V3p6K2Z/0/Lnlbx7whON7XPSL4eo9FkWn0k
wPRvcEAHviMWIQQ2l5ieeWoTdkJs3ynjQ/Cyw4KTEnMi7AvoOt/lmCaIEGfR/DnNQZdQTYrr3lk+
gcBDpll+lyvHV7pKM0e/T1re/ZVoNi78wOxFJsTJOUr1vRZFq9xBMEgiGtku7VmxGQ9c7AQfworD
UJZUTa6SUu5Y5RLa9dWM3JrGHBLEOJxM3jxRwHGbih7qnoqnvBvPDrH/OUhjFpmWaIOyNAKrCCdV
h/wIsKiyIZ2Dvd/YSbpJg3CtmSOGKzi79Xn7u92dM1/1pnRaveENStJvavgG4rweEWLppUb2wqL6
lQSVpvOjHdZxGdu8GkrTk7vfkCPKGd59tpM3kdWQZvBzuO+UuWQLN2F/ccU4NwoJrIJ0aI9y7RwT
r032i6JcbIhNvOtplBvuGrY4U65lLtY4mIsuVXhzMlByts+1cbaMwjdL2TgxRhnxczxCXxAWRXHq
icT1U3W2JPN0eqQFSAUhIYUr0Z0b/FiDFvYoBR6ntN59fudcpFSJALts9ZA8k84LGVNL0LndAYPe
zkCh4D+rpaOgZ1wcG6rzJWjJtFf6l8zx6yLJ+Gtf6wZtO88039cYwuMVppsW/sOVPGTmmeAM+h+a
5yrcpc6N9L/3DccgjC4DEZXXDfvvnXxPAJ0KU/n8VGErm8qsxIHuM2yEv8kzqCKvxhLBKPnkqyqw
eV0rlq+E0qf7sP3TTlT+9sJAeDE6QeAs/VeGAggGsT/uB/7H3BjAr3bjHuBXR59gvRbyczT3IQBv
KQdJVU35GYTyPUZMnTaOhAEuSw59itkigqXYxSg0kifsz6bhm1qj9M1B2w4+ej/TW3GKJOMHtBuj
1HyJBxBBvwU0F65IEk7uv17ccYwMT9daYAblzRFZBBGSNVbu1+JGvVJUbuC0oF0lt5kAmdq6TzmY
OVnCtJsbdw1/Uzuw6i5Z8Gxx6oErN7JDPRWMtqPA9tcwTOQ8YZbZFbmNHoiw8Ta/y2WGTtNxXicm
1afrakbbLTcz5PyEA4kb8BS1qXeMt6z5XWDbkReIKQsPbUgD8m5+ozAShIaqjSmNe2HIqk5FR6dc
CAJFgDdxApoyag2kNWDKdQW1YBouQvwzmHEIWJgPiIIDGQOFV1MyyYR8uaj0fkeOds9pphVyLQ5S
k6iY0JaUwjZx0/FqThM7LgkXXC14tlU3LvmiY6m6iFzSDVdB9j7TwJzj5D64YJj5TAiKlD8X1zbj
4Ws00fCgaGt+zomZYw1quCIPBHff29d4TUDNyyRFpZ0dJ/WwxQDIks/T2nKuP2C4TO7Qx1ETYA1G
lQwXIF2IdDAdPq7zTOfyaFs1mP5atCQNtKxJPItbzmkHsnyg76zdgMsQ4ZoUQ3El04cgSZOp5j9C
a26fYKUv1SDTmy3F8FSyrQPFqZrQEan/3sHB/I8DpZu8JJj6651CCSdxxdfRAWbE1raewFKKe/le
MPWT9QIgeOOdiF8zSZEqLA2J8NT0Hz90nQxtI9I2TO/BxcALavC9o7+1yhuCFwWQzF6UOLt/oeBx
2AbWLiQ50H1PS0WbnRlbAGy3HRWpWZSFL7lVWNteaYDxB51stgEqLcx7cLw6CaM1jRRfgSE0karT
s5+6143Bc7t3lbD8gz1AGOszle2DwUqKx+fIrP4IgagR7+NyXyJ5IUdUpxhnhk+GjNihPE0GSjYi
Krcwy4bL5BZKupw6gFM0N/+nVfAtLS+DvR113LPks10onHbVDglVYROh4+SjgKI57LjRTmMsrExv
cGogGYE3e7vwaMEa5P+bWCxXPcxK22cLKalHpLlAc8HsCtKRrTQDuwue8b9u6KfrDOmdxeskdsJO
bic1z0tZi/Wkn+rplGcJgyUp8uMUtl+IQv8WFaBk4MnI2ycMIJqE0vgIVeP0VZeEA2mBIF7RAjlB
o4TmwS4e0hOY/AogswJM0isQV6NxL6L0EK6ed8ZjztNtoIJeQTzBVblnJwA35o6ZvGTk8PuCAoKZ
cGbb9Ove1rdPRxN/iOv/TG3oJs9j7mwZ8L5yMMRvG8Fwwubju+vXBeFP+RDyNgr6uJUTZm/UuaSm
jBRACUiQ1tlwXJ7I5mNZ1OW4LJwXY7Hwj0cHxkyvaWt/Zwk2yc0PlwICoVXSFGd46OcnYxFF6leq
Irt9EnxmmmlkwTxM69ksw7K0vMcdJ9/DvCSJBppzDI+0AvJ7xOInY6ygA71SAUBVnu5/ocnN6wRh
WBpWWAGQJboA5Ti4WIzC482YVZsilGn7vKycLQoPykezrvZLmAwvkjcIeNE+PF/HjAjW5aWwMd/v
zXXi+DwxKCK0FLiTTodqua0nXTt9zKgiSsncuH2IVXO22QUd/74QgD8LgbDAtz2j1Rb/KQ2FrV1C
oT9G7n2S7o+fX2FqCuCcW9Ibxr0nCn0wXaurXIiB/aRFMUHXKeOO4xxBHypxqLO6red0Palt+EzJ
+axAMGQMaJRVB6LrKDcUYJ0fb0qOIRJbuYFu4+zKv0uxdgFhqE+pSap4fMdHVfWDsgLd812Ps3R9
aMaIHGd1N+FgvCuKBBn1Qw+NqacF64kbMoJZh9LOICrxlcnpyoDVV/kul4dp2GnnHls27ZxHv2ka
Gzn1NnovxTXlnWi0bjra3B97Ze7fSyufWHvwiQDYnCDwKhAFHlmv9RYb3AbruJEii5FXJJ8/uINQ
TsnpTBYklgLNzLi2dPhdnhXikmAYUhVO38zFeSW8d0/Q8XrOWj244FM0eyAcB5qoVvK/FZUh82ty
w5WVc8fM5dwmfiXnVq4WWIZDGH4jOuwRUGGayn5+z+VQqwXsmlRx62wfS2Vh+QUbQMh68TtbBotX
UBsd/FAuLUe2uZHVndjvsW818HR0LwvDQrJV5dpgmjjnLosOpJaleU0bYiRi4/DK51qvFrADgTYI
d7v9ST4C+HRhtcp4IGY6RG6EkeX4MUoatFjEazrZL1yl2cDVTtE0T99BAkdLsmA9b5oo0vhkyRll
geDX9ert1wOyMrSIwTSTGoDaRpYQELj9EWBfXh5vFu0JrRJyrXdtZ+nWoHyZ2CKQ/epFbt4IpB5H
Z/PWM85uWTQ9NX5Q5eFVtn/Xs5tQvtTgqmJsLEF6M7ZiOgdbvNdDXhlzoz95D6TSi1iH4+NnBPDe
kdfAVZQ6MnrDttYjU4IbICkiBNju6dxXS0sWWmnHaDDlytFMkf2h06ZCg639GYKafJL4b4KE7/5K
RBRFMNW507CSgP2px4EYwXv8zPRsfbv9vvwLYRInb2bR8ZCBpZNyaLyJGxJYgBNs0y19JxYfaHEk
4M3I25+3hGJhQP7JMo5LyIa0IYCMQWKjNpuAYsAg122p/RqglJobNA4r9EvvVa58XSV3Jx9kqTOO
mhVfCVJYGFRc0wCNcnlDdUW0JjiGes/6ejAAfNw86VlmOmjDjTUAk4FammveVMqHGcu6vS9Z3a8g
0r77jEee0aetz8RIAYYPhRRtIo/2lEKQBukoy1JU/FSXc4qvnvfLxMadrqEntZ5qDZNIO4VFrshJ
msuUaLxnBTji8oEWW9WmvLz3A/NC4pbam7oF0+MuCDZXkZqHayhe3GszoqpHHDeLqWpph3ArPbsw
qBd1Uzt/LqIf8gFrBbCjpwZLInwYrlvGgzMOozlMLnz1yaLwZhtLtg8ECv39aTtaZpfhbnBs0rnR
f82+SqARvC9XVI2WLRLtR6I/4Sqr8BpZUV5p7zOMvcSBq3NlD2csmGn94IVYOuOQSE1bYylR+WGJ
DVJTIp6z2WfsLZJjxGhVOqvl33FBnR14Wj8Y/VXeQbc6LXVx01drr4DtDCldbQeYtU2txR2jZusO
U8AirvLuOvsCFyPHPEuvts/sQDp9t7YQQloX9ra3cxlX5yuzzkx2xgwz0pacogJaprYHR4DHxmZN
p4erGgnj6EtLA702h3eWmAlHFRM6v772p24cSzga0hv9YlJ9mNPTHaDAHSsFnt/1nOlN9b9Ttvcg
oH/+yRBkOMp6GLCQVvt5dhMOTSWIzDxO1N2jhaO2ZWo3X0vQ5mVqLCP8KOFDoW4JC9SnK4i5zUti
PMyoqTW+pHlTwpM/qtaIY/0jYJqMbDpgEuMGBHWS7l9fk6wEWYUBmQTOvUn6M96UA6Mtv4+gng1Y
mrvtvgAIymRh7EdbwLIdIdd+Zpg3zq0pDUS0oR2oinFfmVF2hDRN5FfNwETaDsA/3V8pAtV9xtB+
8bsSRYsajc//xtzIfaaq7bstTz6ioB8j1aUftykLFBeFAIzv+ZAI827PUIxmx5wBQAx7mtzHi2Ol
zFokt/WDKcQqzsWjYCUt2cRfGMnaZEi+HSGRr6+92lfV/61rRCbCQB6TDBPXXf2f1MpJJ4as3WSf
w39Tz+pKMLt8yMZTt3a+GOi2o55+kdXTMo15BgTAL1weig+2o5V/NiCgVq/BKDi4SWqqt4gOofsZ
ymn5MTuAWNbVtf3sZhTEIxQ1XGEXIIrb8esdmWqp9CTfdbt2L0bzWkVRb3JwO4Mi56XstYUnoMMp
n7nm5KD8OweCgXzaEF/ml3HiD2+KB71AD/IyFRRUDBBRfqsYSKS9K4OnxcJfYHXlwqT82l+n9plY
erbuBQpRBKYMr1ejp03bUCeNKnqCXZSayS80Amvb2WuwewPMP5v6+tJ3eMHIpGlWh/JJcO1ecdmw
PJ3z7lcKVXQQtCHLFaVdXnnhouEmt9iNq6yDcSIGLh51fYtTriLxa0rEC0yp2UQBJOIviR7ikd7j
apOJlHUJTxlZ0dFobDRmxEN1nNaX2DB0i8OITt4UA54ld49lnN1nx3ICcOxovkfvbynYtXjL7BKs
dmmLOFnlINcTR7Y2LFdlFzGFcqSoDhO63Sf7BrW+zSYOkY/I3yZn8z4bGU59Bbdw3OZMNOAvRBfl
xyUQLlUsgUOpfSPfvwo8awzOGZeh+rFW9gTCEr1PUcVGDwQDqV3JX6Y8Dta9wNMFekHGK1uvlPDe
r/2mU8966jF7NTbY3i0T6963j2RQeAdVU90vJgcc8OOdCY24wS9yfSsptrSXOMcSvBlbeB7vhYok
eh4i8jVbK6rPfp44jAd7bPNgJQ7VTxkop6olbdtNn9pxqvcQv5WOQD01lg3lDXzX6pWbvTO0nkda
JAMRREf3Y4fxLwFbB/p0KIbuKx3H9ZgkmDbLGp6/yU8LUYJiOu7f9FAFrA/C3hBlg0Ek9hLYDzpW
lsxVTtIIppQQbrGMuRnb+/Ufrs+kaUWPcHGSLEUFRV/lIcsYX1Te09Z8SiTrZYE2m3yciaZcIs7/
RIEu/lY8hS7nxhloKL9/P//yX8bxjaCWw05FhLXUWc246fV4K3cImdo5kuc3aQtq+tTGxg3PkLSC
M8g4rkZb0tq5D0RNen9W7bB1Q0N1PC+aczi9mINTXzhSc8gn0UWFi7o+IwNL75yV9EaZmXOa2N2V
MqMu9vhcxi3AkFJQ9ZQDGF4BCqfYAApvQyNd/LhMtJZREXlnjP5g+NOO7pQMaqiq3kGsc/rK1Kps
c1kK/Pw0zePeV/BNmwnBa2RDmPw4buCyjgTtuJRIEK1O8kEy6f78eIkn1YDJRnoKhIXF4Y/I3nVQ
XpmayuBFwrc2zKj0lB4EyC+VxXwuEWaO5K+9AnmGdU9/FpRahrkZzoN1ZkSbJlh7IXkIJQNhfFFT
wjYZR6bowjMu93mjHl1WB4srf5YQAExtUpGeKzUH3AzO54EIs0Qea0gTasg5Y7vV+e4QHoF4CNBo
+8hpMY4h3BdRWGiJsCaauZEP9a5FYqSNyFYvyK7kbV8aA3ZjO6Ew6rZ7XpIfEOMOAB4iW4gNtTS/
YytWkH80AJ4gFw7MwDmkioq/PpFCyTAoqqrbd1IWN2z9IVZh8hggexlKCSLMXgfoeAnhCnSE3zUW
F2Cai/QErb66N7EEEOb3AZAVBeOu99KB1hrImvLApfMMeQ7vcZcSzqDIu1kn1bO2/TmqWm5Kpczt
sdyc66NUMVeQXmZ7gPE3GUe7ppT7tKJqu9lFyP2rMx5FTVzWwrR2oSaOC6HP+TBV+yYXfIyMEgSx
1O3/xHIUxJm6Fpo6iHS3Oecps0RzdDh+ZYZfpr1sZKsRAhGqQ2iNNexKjIUOf35jG8B/GjF8VXMj
W/Nwa0/rMBjuQHL1gUnv/RVNIYGWvEUqELLz9QyJiUdFMzkfhXggOynypSP6+Bk6qnHv6sbueE98
Aq6ewt+B18p3Q4N3CG4Gj7BkhmkroOytZ0dfexq1L6JWNk4/FzYvzQymfG33Ovn292RwsO6eqjqo
c2/+OwD0xH297xApgOXUwKGg5zKG/5JhJitXJFG2FjjhkAlBTbTG5baapAEZjPHmcX51yDIukdau
EEscwoldmIQRb4em89PkhiUrrOY5kHY8aHBLMXd399tMSTND76vyruQT59NY6YOsAXBoMW7IofzE
1WrDJMfXW0fvufT1mq0wbW1hOfKMpPcnjwEliPBug+wE+lYRCsYoOwUGvi40gks8DQ1GGAggVl29
vfBkP2SVZQj8qkU8eD/2kxdBH4mcNmcbTY8h1SXhbxFTnvvoDj8CiSUjVYGP36GBlnU9fJr+P5vt
vtENM6p5BlqUoh7qal67NGC3Bl4wDjLoJ5/7Zp6g/Qut3/KEQXGBkA4sX3DWllfPExMecKYLS5Ib
RFXomieHDhWtYIZC0hgKwl+7TcFq/70ch1O33Z0xmhVQ4GCL0c4LoTeXEJgbJEakxFCGAKtcIjbM
7GHXxol0kzUj4rXnu/XWolB833oOUghM38wbzllw/E4cF4Ky/bAB9nrGje2CoQFsADLGQTEkFQEq
KhFZAlAbnY0UkcvR2kMJZ03CFFWpSPhrctz2KgWeH2ITSfKsQptcZ2oqza+DgVY3s5omg/Ehts3U
2HHbYCQKJF6OBb6VNauvVQVjkVRlMDr9VnXx8zF1Tbe7pfx/DOD0v6hYw577Gqm6ej46Md07OwLu
cYtNUs/y3p+UYDs9oPty0kmgBti/ff6hMLEaPWyE0UAVwTB/gpY9xuUY7czTOr0E5qhJtxghFVuN
pz96iUHa59pjyeh9F9SA77R6K8qmPWMu+iv2ipdG1GrRJ5ZamXcJPR5tG2Krc+T6fY8OZTTwVEpj
E/q/xrgSnKLGAh3hm9KKAHfbxiktPFUtv3f2wr/WJ+RiIrprthkl6YNlkq3JXjQ4PEjoi5QKf9cJ
vP6XelWni3mo63byPKSqXK1jssjk8FsLlApPFQ6Gmtgmn0wR9lXuDnU9Pe+Kqbuw/s+5LvAG49eU
AT/n3EXesRnVNOfillfQisjX6dpIi85jrWGFEoeVD4C/EXBZT4pB8hL96pyfIGvv4IelwUz3rhUx
idbRwRV6IEuuiLsYeKPLMM2D/eTSa0ONb+Fp64Weg47TdxKGa1Lwxa1ZEG94ACE4x9fdQWJtYSb1
ziZk2z2xmUaswD/NeBL54balYntKnOfjLhjQFq1vovvuptrwjLRTfBTgDJdVQ0EdAZGgCADKuEqD
5X18EBGPQwN959IVOorUiADCd6aHfePFuxQf/WRlHTh5oWhHHpJxxPmq2USql1NY1kOn5W0X6ghS
EQYzLVHD6/fqnsOWYfeNNeqf46hHNprnBJvgEeuGcbkLIlPN7OT0jqOXW1n3JtlzXJxAU/0oy50X
yijbBdkYYEFcg6h1b4/rJlHOcxsAH5cORd5s3pT+D+aVBolVYR7gISr1neDONVxMGl2hKOARNpnY
a/CADLqTtNs4BTsitXc0h+g1TFZbqukmL7nP7uNRKxPhkpJYBpPw0WwOdEsyZFvQ+FFB0hLmhAP5
BFXnJLB5yRvdpE8HQzUBid39uFoA0pfZxnBY0bYdtzPrPefEnkTh1VWM1xyzw3PWzkkJZvx7pYyM
7VeoAWsh3pmNLp3dodWQx4jLxg/bk8wT8uKQmT4eKE8KinHpuFLyJhO0LTyAKvGfnvOksOb0cY4a
phJdesw39SIFzQRrwPqAZevpWOP1UoldmbYynh94CJ7NsEWbH8Mo11tw2a73kZo+/cLVNtuDYvzl
700AJi5faita3/nr5HWXifngzaPBu0uC9UCkWDsBwI1tGJsmlBdqgs4upRm3jilhAudzO3r/oJt6
pncF7NmCEncdJzRviRMQKmD3QxEvPabjdO+ayxJje2TH+Uw9Ieiy1dXwFXGFKunbNH8KQ5sGcimo
WJbTMTsi0hie9McNzCosI7pJmI0v5mckUe72RDYbNq7hQHTLMFuIShVKdWZf62ao8fRebZ7de1Uz
J99/L5yzaicyLiQRAAlMeH52dt9brFe7SXdMx/B/USQn0FttlnlbBr9xJ60YpNnm83TrnY1ABjgT
jVpXOxsBYY9CZufCQvkCFrotoks+kTAM9do9yTC05XuLTkgnQ1JqRQvviuyOBItMYVKiEyTcRS9x
KklSXddvEp52r4Clyk2L3MkMf970Xuicd5yFaCBK2kcV3NPoiQpHDU74FXG9WJ3T+9pWBFZz70KC
RkIupl+2CbztDus94c+P/cfwSlvPIgvIL/Mc1V1w1h8kPKzUJE0fEtDaRvbzs+UqgcvbysDcYmRZ
1u3lR2EUvVS2Eh+94KzQoPz081pELgMcxLf9BapRCXoJLn9fl/vWCk/1rFywcjkOU4QxukmnHJiy
WoRLi6PTnykSyU3eUiJVYdFRds3s2Wt3kFpA/lPdDwAXeg4+/YPEu/F1W1e0Ir9B5t6OKl9MSNN2
SBasMgUHmZGWqjz+7HKnKhrSIeDYWdh3Pc+avjO/Y9xl+qO2OXocbOhNagGiSDvgFZ+2ub8R5XY0
n0UycCVfwoorerDRHeuJ+DW4jvWrkxcgK1fcth2JRXGMSJp3zHu2JaEZ1p0fUCKoSSRQww9xpqBj
ggLHuVCQtx1f8o0Er4P+kjGYPabcz5HQ5HT6CyOMjWW9lhNur2OSNu4t3Lo3990qmmqBdrdyzPFY
x6XPfBS2zL3SpKGiKg9+krj68da4Uu2FMg09xHWf7hAk+mPd9doGMP1T02a1gMfIZmosVG8UNiQB
/975SaH7Y5/aVA+auSwLxVDL+FWZDq6c8uvNDACBAqdM3m7UNNNLni+OQ8lPudy24mLRZM5ZmHpI
6DaZPHSYbm93J9N3I+PZOZ5+zlt8CHeRmzA7VmuoHJW72hsL8F+oPlOEalPiQFcNceYSzcfqJvHE
xR+yPmkG3FhrbwL/00Tkdut2qlvcDRndU5u+jkYUoWKMbr8HjPRlY4NnOo4xRLNVVRq6zkbojwd6
t7fTYJysgdSdGj49uczyjp2PdGZJ/PRWGannoFWj9RRo4pjqFBroiNrD1Xe1+9rRLvhGr3xjO5nM
Pmfr6ro1NzvDDFL7iLkOtbPu6zLAyg/MPewUI10h1FPd6aESUObGI5efV4JuktoBkfYyuBkIEMUG
KgM1Xuu/IZwcwewRzQKgWcXEDUeZbMkCg9m4UyOSssUGSyOZGkwrp7mScKrBXfxGmXmXOPKoXuev
2E1Hoqw/vLJ73EGHBlO4zAx7BISC4jN3rQZts3Yz09Di3zucdq1otxMfrc+hlI16sbIp5A+frEe6
DTChj/clKr21MOSMkTke86IL6hHjaq4342KO5hdxnrB5ZfEtTGotq2GM662Th6bjQLYfaKhIs7Tu
n+4m2BIiQyRirj191MCMQNqnXfq07KKyXUpz5Plc3TmdtdMoL8NqLwbqR2F02GVbu0E+vJRoMUie
f3MpPOw8ThVJl/R6HGqh1emj9AqiwihHo6ZUvHvTbXfzjFAFGI6xgFLk0OekUACcXY2s8QL4kReZ
FIX7YMUaYrAPE5gHH1teta2YITAFfz99njOy9GIyW1msapzrUOw/8+PLc4DG8mICPTtpChn5gnTr
2XzA35YTj6gMthLEdPaiy/gf4Yum6iw3HlO4aYlPulpWLEEJtQJOQRGOzngqGpYiJDlBM2RkwhLl
f9n8AcksoqyCapEJLFBPIyQMRrTrl7wRfSZJOKGb9kHRDxhPtya0OObnLD5+dTbq7i/RD0qmxEDk
drSi5lAQkZIrxgKtParOKagnaY1YHL3ZqMX66B8eJJNxgkN9ockL7JR0GQ8yJM3wtCOnKDxNWO1S
MN4P+DOQEF90iM4ynrHRYlEgsk1/I7SRGqkIyD69BZ5yiX9TResszMKnIr/AucqaXb1T/i3lLc7r
eNa4wOFG6As3mLtuVopYgy4hFJ7MV5zg9MnyTL/HFNDRH3fY+dllwCkT56RF5MfDO6lJv+J/Klps
GrjXmjr7+ezhqwApLLfie7Z/RpOSgDJC9Rts2sXciI0WoOiKZ7LFVltpQUM6nbcElhUKbSZVEfGu
/d4PE1odRwOD0jx4Xlw0+EFTGitq0kbq+hY3mVQu9nEKbDe0N49p8fF2o0kG8yOYkJuM3V6oeAIC
E153PxfudB9mjU2O0i7MjbDwO0mBGW8qqeY7SgB0LZyGtT3t0BHNNlumowWOQIj2V7Okz4Q0ypgP
G7qGZx5tYUtfNJ2FmSBWx1dWiKjOczyQqm70yPBLX9+267c0nSbm/KWMB7T4h4YRE1PEnlNmcqlJ
WXSaFsK5cUxLLv1VJ0wjq6L9Elt950GqomzizqB6ENRqarxVJUJQH8Knfmmn3bDHbTZlvD+8I6TD
MBdC3EptpcL+WZIeEZeN4UtN3HliZUX3P72INKMZYZFNiFwaHEhs41n4xTKghiXlwvXXUdgmGAEr
+V85rOZulZ+BUar3W2KbaIL9xvtyvJgx+PwTBdNW9xT5Awn2JCpxgsrjP82ddSE+oIhbuAcsUmmm
QtEU0cId8mbtTl+OqsQKQO0AtTxPSdCpTl8E+vEbJW3FgpgOZNcPVzN4CtzjGtk7SbSnn2iAxfY9
7Eymb91jWZWXN7E0XWBAchLzk2mOa7usKzONwGtCmvzFOATfFWbYiMOLDovzx4VrmVCV0wKh2yxh
LAxHtUCUHwWFCsBp3n1318eUCxTLqytzNydER2v9lR86mVzJEYx2Th/uTo6iQMLoWUwPOQO7mPCp
BDR5Ms1JEfERbj26HwXh9T1R4yEJrwwvPJRlT19tO2LK1MTGbsAolO2hzFIH1p408BKqdtoKljEj
j/xys/yFXrQYyVUkIT3W7XGdaIrnoaFV7MUMO3uweJXXngyfOgaFbP0WTfn+qyjEGYn+kP09Ycq4
kXIs1jevP/qR3p1/2K8o1mRXtAl3KgVh2W2vcJvvsRFpbJ8C6BNu/XAreBrhYIcRFNqyvqQ8Zktr
AW/eJswU6RNgYWP9YTTtkjUdiMCFs73gFNGt1xyI7VP1ANHu/VGE2XbWDIqze+MNeGERjljlnX8s
K2wF/6R6Gh2K3jx0gpnY2EnZ4rJT/YHo7Ls7Os48WZjEOLnZErQZdAOytrdmfwzX+HABQNcx9nF1
aS8IwnV4lG8K6KWwUpirLzEmGwu6ZakodhqggWmgB2uwPJn6a2fVaPhC7Z2baIr/9F7TyWFm3BrJ
sGoOU77z4cAwe0ItMg0f7sUkRGnbi6iPLdQVYcmUS5CoJ3hwHQkCr1k8+NUwhJlbAAxf7mhKu7rb
ZIc4SNZbqOixZUirAkeoiD+NkHsDFTf914ZvCiNMkq9j6nKJKfndcdi++Yelic2mCSR824Apw55x
EJX2rSh9YrdGG80qgx6P7y2m64UKDjtJZ8Yv8hiak57OYrnYmQkyC9S2YWNc5oWeMHyJrQpjEGzQ
o7gIhofYkQihJoX7v4NxZPxPkOAbhJn9bHte3Vhr1t3SYeJhNItwRVjss7VqKIr2lBD6xvPo7dlu
xjhs85IpYnYVEVnU2bKocfEpXBh44pQv8W6U2XNE62TO4nssHK0i862XevJ+ASadNB2JqkhG20nx
wzuU9vJ2sPyLUKqswMS9TUb5iqdE6uEot7fdm0CHd4JQK+u5yzXeDEjWSJ5/Wpme8+T6KiZlyawp
sxv1XiBKfisTfNgtTQq7WcmE1fi0u0z4SA0HxNTMUuQVPrjPwb8bUZpu/pi/02LI91rauGagFAFr
nwCNWOc2JSrd+y2jYE4CHdlE8iOWy6IuSxXp1eI1I+uL1VucDAHzsL2geuke0AoHUIZAYzmvrgFs
a4W0XP2R6jyBdd0TSI68PbfAdAK5TJmqZNL6nBvML0ASEKSG1aAu88Kmvsuo2Lvqn3ihJvUMbtty
7BsnxDsX3EOairNKO3Oyz4wj/n9+p+r3YVQzcaXyeBKEJYbOfwH65b7al2i3xv4OE6j/9xFZ8sAV
cDVE3oeIArM3mqWS3yNMgMH1mYNadlGIcsIxhmXZXxVX4jgBnSNcwXbq1D8VxWgo51qcNkQF6UbY
qnYWpyM0QausGvH50A3Z7TGSx3rzpt/Ffed27bM7eM79c3LBIVv3z6hs4CCEg5Uu+DZdoadwnk15
TTcIhMPUaBdzchEzhO7k5ZkngfwMluNI1jAWt65IrnbN0iQvaynLh09m+tzK6FD46+ACMSIS9jy+
6gPEsPsA4SVMLqQGhnrYLucbRp9gZKlGXKvsZ0YI5xgSX+YG7xzYX1NLXN4tBDEIw6ZNGzfENy4p
7oRWwFjwbZMQmWtmzlTQvn7JLx/EHf81vg+C1C6Bg7uWzvcNPGs6u4mBAxkXLBFK8jHXq6VK4+99
ciTcgg6mhG/KDDSYXNCMSdGL6FAGYKoptYRqX9crDr/xpJReLMNGNw4iBmuCXM+t1eKQ2jN6Qima
pHNvBbrlEl3GihlLJHqCBoDfI8EDz0YEUvAgOVoDc9UYJpDSM6lU7hsryCrBcbi6W2Plj5BjGwXn
2bE92KGpSKyFO8HFJbkVJR3+DU/EjhA/1979D2IQjNFlX/dhJwzx+qq9XsYulXhk2ZfLd+8o9Dcz
8YBmyh+Qc6xl01GvfIQQOIzkYzOxO2H8sYszZSidU7sUb5j2QpFc+wJfyab3gDGeYEt8qnMd1KbR
LgTQaNwDrmmg4ZCcd8j9ZNHObnx397vkWnWMeCRNdSPetPM9ukjaERNz8zqiH3sLUviTf1CkndgZ
P+JJj9ysAQmw8fpNcovk0yHg89n7283h/dBwzseq6c5sV7jJInpHv8ZhVWq159GgcZiiX43/gGMI
Hha3Lg0PqznnbIs2OQm0IFJWUe/tfFgfdenGlET9mm5lMGzlc760+DcNfQ0pF5WnjiYO1dBzre4W
/a6U3vO/BndNmXzutaMoCe6lJxvs73S8xGT5sjQ8rwZ9+lIavMr7x0nMcu4ngrLgufKAFaVnntTz
uifPQQpcNcZSVMFiO/+LRMw538pqPdzW7enNDhmbL+qJBGjFIbJTwuCMl+FdEG4rUTovYxkeHvEv
lCND2uF2d2YGKoW0lQ7+7gWLCbz67EPX6X/eEvqDWWwkyehHZQdmeHqBFH7qBgmU54nSSOo2u5Br
JzIbJPHSIh1B/itWyNGhLEIp0K6i+XS6CRWXL3R4o8gcgU2AJv2TH/7f38dJDrz+wEJh19o0EPi9
RKBMC+w98LnSJlYCu6dbtgwxA46tnz2SZFbhYSfu0lT6JUab3H8rtJCNnJLDNa9uPof7OvgQjP8L
tPyOXPR5FSJqMPz5wp6Ohb57szFInB5cBf4l4bvOJV/WqgpuUZUG8huIuhYGSWaIHGKCYy3d+Eql
g35Svk7uREM81lbhMlAXEtEtPt1N1/JKTZh8IfhlMDR4jEaYLkcK1E6ZNqBvTrmkGoGnunvW+wI9
6al1aj4j6kkI8kzAxcgP0SZUfB/J0CjNjFJxwAtXuXZnGDEczYmHNyidMfPWe7nXk9mZEMnnLK+/
zJFyCWcwauqd5yDIGiPBONQVFOOrNU1DpxzdvFgaOQVcI6sUXOyK0EdLnBmT02mQO1+qKDNqAWTU
DK414wd/StS/RlDcUx2ylGDGo/YaWkbscJZMiyvG6am89trqQumEdvHDwMtP/c5/nSHZ2JhMuML/
xqjRAUrVbJEygoo+9gRwpeb+L+56MigQP+8P3eWX+dcWLpokWpEtXzZg0+/QXggyqIoeKM7Rko77
EPrLDxqGqhm9TpaASOfiM2RvSJ7cAxk4H9+kWt6ozqolznQ7xO9a/nDTMGlOu73pUBdsqVvrvpTR
e98V2zErzhEThETY3e+RqGfUoDV7zykGRx3vee115Uqzuy5k2BiBIK4yE0z39sEtFD6H0Qrvzkxd
UqGx4NU4AdZDXKy6hGeaqH7GLltNzQEWxa/etkzr1tyk8ne1+hJySyAtt0frjtq2fEQ1+iKnzQFd
gYspje5HoVs6HPakix0oP2wfBj9MDBMbiS533mBVZFjyB5Ab1XOKredLAL39ZTtYnk/uYU+W6d2C
MohxqsIH/WVLGewP9/GsRDk5OqjWm7P7MCXcHO82FKv4t+CuCoPgh6a4D+9eFRqSQSWRm6zgfd1b
45YvQ88zZAYzIKLJA0gSE2IJk0b1qFq6Pz55tIZANlSxbdndgceAeHlVTuNcdlJH8/onLQDTKc43
aXKFC3Ffl/m8CZeD9S8PNpCL8Ts9r03Qlk4Gnws7jylIihtcKzkgxhVA/jnLzxj/BdwZOU4mOBEN
dnaiXiWkkNHlFHSB5Bx7SBZryJ9lihriv3gjpCSaZRC6BAZdGP6D/Q9HiRlv3fhP8ma60G8RMnAi
Es8D/g+NbUxJfQGydUeIFYqQdFtkw4xuXTsH8A5mEPl/WcswpwPyrp1WcaGgmtHMAvfQjBbGBn3M
UHLUAzatqUIcABRFRuV1vHoqsM1nL9JOhrfrW9Tr/q51uh5VeHPB6CfqnMhzVdmuOgXjZSWszsOs
iaM1Geo6e3wcQC/Bd8NPVltwJgYqwx1ag3hCdwA7tFgRAZXAo1opJoamEWu6i9GX7HmSyLEE99cX
gs89q/rL7nTC3khZIrOJ6CVR8L35xMB4ISv9PAuu6LU8w2/dU9HEfMnfJDlMhCsrZ5d5EVo1MuXx
ZA06WWtXPSlx3Y4rhOPA3twlIVSu79udLkGY8fayR2G4nWY41itH6QYgkfhW4poIpS20KocqZV2y
uz+1WXiwqIXbmTzLA9hRWBITtFeMSQVJy6Mr4jZ7SdiEOAgObqhhDv1dtwgsqDZRYD7zKGsiP4GQ
Ffd5MAu7wYzw/d3dOGKh6CcMJ0LQnAHcczUpIR0NY9g/FbabAKvSD34rAeD4gFKY2uem/TsmNHIV
TM0H+s7CkUq2/pdnJLD2Tae075oj9uSUsYFKoIuL540ODsEED4SXcorVfp1N6h2VKZGFVSxLjwCA
yADR+aNeZYklqYkgULauRs5rnyDTKpDg7Ts3CmSJ8tyFYFHitmTHNapZdKkaWeVNVtTpADczv9HY
7LwWAqbeg6eomYxNMeviAHCMhh2ey6sRdNCB+j/VSlozpCaiZltFX6zH/kyJWnuFajsyC7c5WTXO
Yk4sbq/szMwfVK7ZB0biHtUf8XjkBBlEJV1VmvHGXZ+0ZmGiHkv9E6JyKW2MnFWNy9xn+Yty89xU
HHtfUNO6X/ImPz5kso6LEq4LlIzFHyBaN+3lY3qmenhD/ETpnIwA1nV+D0YDn7/7il/kCEP4Fmfd
nrlbCnnfoTfVnmoE+pJUuI/PIZJeRKHxqXNNZRYdFgrZc1+1xfZg899NVEkzeyXGId+nmVeTFQIF
iXY0XXjC9jgd4mzbdtdLd5hKiehmMG6ZCSwaIS4/awV2CQazWMNMPgJIeL0Ig9XpAITlJSBMH351
cs0TK8jY6vBOLEVdsNg22+QN9UaVFMslqDdSNtRb3/Cl2QEkRZoG75W4jll5xndDqqglwk3ReJmW
T0iqPzOBilh+g1Mm8IZIXjc6nEWJBAgciBePaP0y76VV5YNXpcshfri3F3/8wEmwWHBmAm9ycWZV
30C68XWnu4+yrLZJewJuqKGwm1N+hvtN0ujjf47hSa1HI8M16L7DktTRGRpGsSnqv/Sb6TeBzNK/
KYb03cUXwsV3K1HjrK+A5QHAiuB+divTBh/iN/3+pt7Y88Klc74sDLrvc9k1TeOhAOIjqjdK4Bsc
nT86OhYkklyVzzzN1CgzuCNxk70gQt00jiWHM5qpXSxqcm18JEJsfElQHA8swEtB/30rWLMkn8b0
HKavSHPPlZKlcF0H3I4h19bFvBMa8ZxeHFmz1uOy4USy9NMrUufTtbUU3eAd6Y93gYNYfEBGZtgo
Vu2ASV2FwaIfjrKdPDwtAXop8+c+PpSmoEOJ0PSnVA5bi78E8V1v1HBkFIO/BPViH2RQPH/yb/qZ
ve9GYTWzMMcdGjm6mdH9yDtwPzQjaGJxLgp6jQSOxUjTwMa31tR/uKmhwaw8CDjg5wwSDhjmVGBb
RQ37Qy58D/janMgw+6hrzfLZS4YIhjCJiOqgF3qQkMpszKVQXxVRTNjkFTOVNoovT/sZiUOsIy8A
nMkOpqcAWlDyku14XAasjwIXAm2p5CLSX2Enc6Kc2B/TbYZxQfqxWPU2emWre5mM+IRwfegmn71i
3dLwDxEOtlPKODUVxZtHVtJDWqh1av5OgfOUFiVieXVZ5/k42HCyT0Dip3Jhv5WMdxclImsFk66c
fuvv4nF81c7YZ9hKNNjYmCcjTWwmykzAtaNOW5qwh5t5gxr9Kh2+Rf2aKkfsc5FfWQ9Tm5/UDiXD
eZVYt2QhyTYVuJBxDFqLEj1LuL9h2cWHjyO79iXhv4M88YnaFrkHAx7TWFQ4OvH7ySl2Ll/UDEg2
N7LTqXaKODvZ/g2JDsAgCPttK9a2vSHxxqPL4rK/4gPpsmogGc32RdCT0UjiubGABVdvqAPidNqj
zxVD36ZdRYx+8rqhY4XoOeULTMVK1C+V4Vz6yXFS/+D0+QiWbNMQl27dhbe09DPaC9cgmuPCaJ3S
tk24ihrRnzPztflnws4NH2cN0dK8BaFAM//NyxPGVUxH6LG4ec2bRoKWCWVO35s5wOhmbaXkYVmX
0Bqb/xuHburA21aXrcK/LCLE0jeOvqkzQE4dbVpuOQxsTGyWmlUL4raqduIXsZDn686wPWic9Jd9
bmm4UW+51fNxrAIPJDehvMjPggSd1V04EUNYo973NQ1TePKUrKTJfumlkt/XE8PvdAVLpAKJIeCH
kJKZHvQJdljNID0DYr58SiVDQlooFGOItMc6Yons9N8pLhJ1AelcmQsyljBgF2kYz+9Qy2EeGtzE
NyEf7xgtWPvh/od7qmV5DEV6PMvNHMG5I13/7W9G3DG2vFrooYbvj9U5iJBPOHyXtnlep0lWqitH
jsAinfghdK1TzxH7jNVEapMLIQWQqwYl66A/8iXVS3X0HVcIeeOXlKHODq6ayM00whMIFM0JUZ2q
f0oVtEijOis0Ny7mLW9jehX3x+bsfz3CEha1DZoG0jMXBpHZ99AFpxTeJtxlZ2hj3w5BFnAZnzJs
ZrmYOk1cEthC3il8px1W9CJcGstOhVOvdct/qk8bZeRic7RX1/76B1nzTntPSIhT0nfgcB52aR8c
+57Xihcx/VU2zt7vNBDnGBmEq3m7CUyfDVqbxBpVqu2JKmj/xq+yl0nii0qzBiXeVKbogdbeLRWy
XH6SamYUbsIs3akeLWbnztsvznV0SEjQH3vVK1FctCsu7aeic0Z+VZT4LQmCEiDeRp8ABVmL7Dvy
tUG+FVkBepN+t+iz97KB2rwfn0T9YFYOjW6qqYMpoSBWMyzirmys7PKgS5dHGxZlqVrBgiFiSofz
Nz5UlwRrp6LhYioT7r4wTbLZogSAgWoGcRDP5YNhPN5D/Z7QP9kh32kmCGIVP6WqYd8nEkvjc8V0
DgK/YP3ynx9ia1F+XlUbDX5GxtpYtFvRt4t9Ats7bMArTvqVjW1vygzOTDCVnSAaUt25PLfDfVb5
xcy0R4PJoxO0L6/TQfpn8+BuDzgMhnpBKy/05ZTbn0mNAnd4RdXVyC8s7rDy+FtNM/sZy/gnBy3X
1o14B5qObjO+J4Z/Nn1V1vgByXeVS8XvOCsTVMCJT3BxbXWdlBb5MTaeMks2qZVSWoUfnbar7KTD
zfyKFsJoo325ObT75nvzrk0oXLzngVSUgu6c3tPsL5K1pijY7y2C5jg+L2m46kaDKN0uL3uyN2W4
LBvxqHw1tkP3kU6FascG5vv+dby2DqacKy62UMeYuuJ17KL5LL24EJVQZ2slcyko8C0GWtFd2JnQ
TgAeNyY6UzrKLO0vCE6aZVKcfg0AsAIwGYO9XI2mQvY7lP7zjuGyE/t2z8Yf+tKIPWs04mOwtGsf
Q27O6tdHPrNtMASrwayL98e172dd+s3vw8sg+5o25wism4rLuaf8qgsvLw+Q3DWi2IscUe4AdDCM
5YHwOnxLRQfKtJF00hDtm33dZ+jgYLOwWtVh0QIKWvZHiPKeKcJKBypd5xrwV5QBo4vx22vnnIzX
1fr8+vri+ZvFLKimf1FHKGsumKh3WuTCGirdy8vUeTLQPr3wsu3u2tpv+7amh8cUEuXuN0It6ozg
iWLCtaCY6OQ0HCPzdd8Rwwz5VRzAsr3EhjjGpMq6mWwyzpjulwAyUVRh/Tk+kJnBbjf5tDd24jbM
dXycTKm1KnAgyYzJty/YfxrQTK+m7vZuEBR+EzSyg2LTvm00xLnhK2av56SqMzUWfsR0ymBRWvSG
fVBFy5vn4tBiPXOsj8AfuWAnK3Rrktvm5/vvhkGvKZrAN1piGZYbml+zNskRD8UUeHsnZnJ9QXU2
hyCT+Z2K4+vImOy3vLN5KaUkRVEUbDmD/FayEowogymL9oxnMuf4XrRFoagXV1HdNWETSAuhckn/
4RfAq9anuGhuP2XtLzOkA7XxDU4WL++PpqbKXfwgBgHQP5qCCUKxYmdhUMcjjgp9uQEo/eNuTPch
g1Cjxpnpb3KGFnvGaA8fyV0NDPJxdoTMnSrw2xzQi7IXoBmyp9EvebVZlGyijduLQBEv4xq6OTi8
WsFeLJT8zNz3rbe6p2zjjVDvFvHELDFF4IoCue0/VSr8mlL5UQ4UW4Cg4Tbd8v75oCtwCXCM7nty
PXvyzw1WCStsrJBlcakqf+uQLdBgX/GjiMl34HWpqAhFfQxf7FbnRJxbBe1sozp94Dmex69VI8Rc
CfiDC9HX3KDUYYq6Xy0LzvEbhq8EMeIalJaVnN5uznLYT8e9Uz9xAFujltAJrVwmaRCVACzt09iE
g1AAXo4I4e+mSVD8v8z+uflrI6lzCWE6FvgsA8eNqY/BJ/D57zebEG/+Cpr15fkHUr6Pe4/30fyG
2RcoZFMsLAA7mcn7pHy2Ag1z59XB7LkGZUANEEW9SbzzVUqcDCApy1Gv3LeWeNOMXSBBQ5DiOfRA
+6Dr440xf1N5qbeT3vNc/rSZzNy0L2e6TbPW81JMn8vPoAWfxl9fOpMzo4vhqrdVrRdqFT7kHxzb
17rQuYJwns2371l57xsepkKjUTdZzHx8xYANTEU+tBA84+QZiAT1SbJp+JANhJWY2TtfNlG36ZE5
sXiBEMxAZ+b+/ZLfT5TuZBdX1L6kEkbao/mxI3kMZFpYKm7zcniFUmgMj9QxAwU3PcUOljZOq5QN
z6sMjLwTetL0W0tL6vpYOeqGKYsWGUsOrTOr0BmSZHq7W0s5zh6WPBu7tAQXFL6eD13qaPv30kcW
adETK1gS8pg8/tUvP3qkRi4663ryenCIt+G6RxDd4EibxaiKiB3nBi1Kx/2EJmiHGEbo28n1U+gT
TBUTGhm/ALzSpNWXwcY5fZBDw3y3ZfdlaN6v7aNpaN+OyO523Cf5oQqzQqNDhyDj1+zDg/PDVgF3
M+h/KL8kw56HF7UUXIOxBRvfplItLXNInZdoimScjvkGgVHlgSh2o5okBjuirttDPrjFZtyicMk9
RY2eRIFIDHOnTI4hUwDZG77AaGEzNjggErSxVQ5CvU+hUu4xKphU22smRXLMW9tgT8vLcwadQcZo
DOqIRKkElaqAq3nJEWGSpDqDL9XIkPz8c8hEVM0IVwPEiSvksk6mpGQ5W05liTVQVjmPY/JewUB4
8qCmuVhPDOr34cZ2xDzI9dc4aS33JLg6MF8AEv+A1swI3a6B18CLCegcE5kAbjb48wO75/dHQ1d/
sibDtMULNZm796a18Qf3v57A4xtPvTwiFgi8PfH763ZV/e8ctfrS3Kh8giRknJrGnzx9Lsoktk6Z
2BO2XGVxw1WRErcNkR0m0kauE7bM+Niw3GeBMi8NzoTtgzTjjSW0WTc5awrFQ6xn/vNIFmQslWwf
6gJO+X1M9xdaeiTWWbCgPzDabSjoyfm0qFuyWiNHbontEsz+ZLx1hHQs6DqZQ4S10+CeeQa1SNPt
p87IPyTBmhgMHj/KqVmtE+nEFbFcmdlBRuiog+nn1d3F2XJdKJLPbbJk+ofD0yOt3qRDLHLV0dNN
HIUL6GreYjPQtFBtFi+yBmUWPfDtWIVZoxGlYHoIFmxUyTzkqa/RCMhP1qvzy9UaaVpsJI6GUxEO
ioWY1o5y9wsE2PLpUCB8lar5Tg2sLJ4I04OO9JsRW5yIV3wFTRqQQ/hCRA22T9LZp5Sh75X6c2+B
QFvXoSf4o6aILE8a8TQOxM4jETgwW06Dvz1sfuQRqmyslWmRZh/D7PPtspy2Gt+I9rcCzdYsiJBb
h4SD3t4dTBvY6+EMgGTJ0kyAz0i8ZJrKYzE8dJ9i72JYyroPJ/zE3Hk3R6Qvpx3nLnRZ0v6000DE
nZ24Upy1vrZwRW0z+RmeAFijDZn/VSHodAQu+2YDfSS+oEFLC+ZDCwhsx5ZHaSsJBxPAXYDAucPr
s+dVUx49ns7FG0nz77fB6PCmm7Vrw4RGqJ6AKs+HuykxuKjzzRcWgN1pGyDKcxj8ZRBGmK4oSXK5
9p2Z3BjTrt9L6VhfCaZL7L+dS9NcY8z7YOKWtR66x2GzTK85URzc+xn0MHVCa9n+9OR2E+FCwLq+
gGJ5k7XlnO3w6j9ErCOPO9quQXvbUc9Cjc3igyvd/O/37qqz7qOCFxbLpUQ6xPdSv571F6ADqCPI
NdWw1xmlra0mJtb86gwTAGrRcT26J74EjbOdxbEVFrT0pOdWX5Prt7Sp+c+TuX1OIRHn/TYhvdzl
WU6Ea/gC5HKOFKhi6PZPU79hQ5TPTNWZ78QnbgANEg0bY+SahXUA8fnhhhKMcCHEoxoS+b/ONclJ
10NVTpCQw2cPyk3CSpAMLysk1yBY2tEFRUqub5+tPkVkySN7SWZjW+K2v7eKHo4iDU2cYPfEdVjR
ElqjmG+xZdygUAYqTJ59ti31Mk9MsxkVSfaH+0Q1+o3NTPzyNWTDwNEI9NXGDt2ak5ElhQKzmZ4d
joISq09Ki5LcSY6CUxFfJ/wl6y7V2RMRtiKpXEOsBPq0Q2sJF6TKD8+5kgirlxvk38CKqmOH+Fzp
yAm+SjLfahekQdvsw7U5iRP+LRLrGiAkwVNKRJj4nFwdMRc3zBbdvWO/qIs8h25FhZ7EMTAFRQtO
no6qfZIRtRsRaLupLp4Hx0pu88E9NaXpdo2t/NH7UmBxThJAnVJtDIi0vIRGFN7frSzHC5x7ix/L
7Pns3hhF6/cOEJ/8aflPMM8GiAHCBTMoNa6SfIBR3tRrpStazr8jxckLup9BgA9aqqY7CGSH7EUr
AZ6LjoRyR82iKwyWcLJCks1Bt7PP3qlpSJ8B+0lkSTpIBQUVtiwql5pDww3+MiNCNKK4EiDxvjjy
n6iMAY9c/V6OH6O1pK4Hld+rPbgk6iUVDLM5JX3EJy9I21ysMVVYpz5PBhdFZlcmKkeKpdkFTI+Y
3tf9K3Ujh4jOV0Qt7BcTqTfXVAMG3dHAFPakj2DNywlNNp/LV3kFmrRv1n+8cLkXboylKco2Grz6
TMPPeBvq5vwr+a0ObWarOy8Ia6mBXBppSjjHhaSHGmv/FCs9ofdgRa013wEuRjKwgZrXFrtu5hSi
/TvGuK8lalw4UuGabYmVTIWu5rpvocUJeDlMJVE+jrxceCTX1asHdhTcr56n/qaO+Th95ilmw9J2
ekiz3SqnaRvCKt7KAuF0s4vV2fJXN63UfACkgiax7xPzkj3ts2IlTA2eFXXfBLBOETBsvgQXVZlN
+gQ2fiiKOYk1588w7T+O0hkccnYjutNVPkgcFSRYFcMEp9/bf4S68aBkIZcFCSFcV9yx8XkbLxRV
N7FIFzGJBZ3clrCTbZ8jYkK6ugB2CAQPI37zMS4RzbTBsqMh0eZvF8fZJf2XQLrCGAEgrGFuzU/Y
2AvRnmOJEuLaXrO7M9lpEOl8O6SBpqp9ASU4mPdHf+8NMezFsk+JEUdsmYzD9SHsiiAqt96koJ7Y
bRQBctzjRn62NV8LN8obpUx6bGDyMJdmpD1cKOw8jBFtGv9cKI0x+ECwIKK/t4a1FrtP1tZeh0PS
VCDjovU11zSWoXExDImnVCPa/osyjwn7JPX6mx4S3G4rT0jExQquCh6o9wiY6tV6Og9mJI/vmVpL
ixPqzzG+lWvEAAf2l+veldQGLZxyfcdchRygJGzpoICBPcEEd8+l36ikaX8Gj20stpeBHUTxvsxo
ISsLYdlwqPyeJaTjVOeDQ+6KzVKru7k+YHZP3igzZ029s62n5ttYyNb1v3sCf+fOdUnZ4OHaQFPt
b5WJGYORM7peNXLMSzF8T0wemOUyvVubxeN7JMV7RKvjXhgU4DVadszY9inynTL4WCYmbdrZFUHx
31cMBi3ktmSIUUyhHY0RNC7n1BknG5GuPpAxwjnhhOWcMgEZW3V4RwkcVTYyOwcfK6PJ59vs3Dfp
Faq2EHLF8n2+SQ3a4ELlSYIxWid3XPAG4S/oZxo/8EBveDoUxacUQlTtTuYlSe9inBODtiMh96aF
kz+0l3WfVqmKd3DV+Yh4oN941O+r9AdBdsRgdHptkwGqxHCE0RRzVd0dbr6a4mAC4NJWLtbVxel7
ltgAMhnKRZENGLqIVhCsE//GehQYlEG9U0Z4mfRMvK5P02JZu83r4vhzH0M+1fmL/gmP+rvrHbPg
bbKdoosKQ00VdfeJtXKVXdbGmfB+8OiCBEZ9ToouLlyz5hnqWkKLbA5cRobeepHbqm4lU8itzLFo
7MEtJ/f1LvIX3IyS3psaL8lANpkziI37gJrT+fwJ+HJkhQtlMqNyEvxdYep64lHXgpv6VzMK0of0
JUtJLa4Tl0mDI06SojUgDN+fkaWKHTJ+JEjXS5rx9rn3yxwOUjAOoXqkdW/QBnlvQRRtEkZemZCz
wVhkcSC0TZWbsElEHHTvgqcuY32vjwggl0OLWAZRjUg7dk+9UI0zbhd7wFbziweaXPaxYIOXo83Z
zIZqvKGn9UIDjQTy4w9cKwhuSxoamn8MrbVTMhTbwxdN09DM/vFNgKR9wkN3Scpfp0W8AnmzcKx2
vc1Ft5SFqkWa/yiihz2Sbz0bRxOdZDNZ4Aczj+C82O/M8CkxGrjcD/mUdIoWIX3oDFYcwwqpNCuR
a8h3oPi4sb7EXkpOAPmkmm/9xrFqYx+bpJuYBeZjYtt9FGgWgSLLewPQ2dc4pVlxqvtPKo50c60B
QVQptPl++t3/zVMWuggkxFXE6jBJzXTJy1b1GTnbH9jlOuopF608529Kf3Yw7vjCrONT8o/YietF
YYhuxwGD8/R/C+7+cc4TEaixsWzu1xMacB4BH+sn2AFxs+HAGV+pMGN4wVupfZaX3S9gm9KzQ+lN
sA3reBEnMNxX+WDUIP2fs3bKSiXvTghq5bXqIUx14b2cy+TrWDtASGOkvBGkaMqucsKFH03cBI0l
Er1eoSXaQLgclwHHobIDQoLWDUkQtyfdDGCfJRiV2CXjRfV/vjhlixfvb+10VYkms1DPAgShwZvs
1D/74yXRalrvDkWn5Z3utQk4WRw0AmmJMoq7sRbvzqNadVIW/dcnwE5iWksrF9C+2J6qY5A1CXH9
yFFLuWXlYj80DzSd4qI3yn0fI5hnbd1/r8sNqtPFgFvAw/CPc2AURG1HBafP9zyq06Zcb3CK7FZ4
b8Hooamy7CVXUGF+2Mz9KTfrgIHR/GgMeM/W5zi8QsRY2SC8RGvbuE7rEc0S+aJ8gvTU/YkvJp9+
BCRVgNp4oWETKkSaJIsvDyPOfNvz2Hpi+bzQ/MsTHULcgbASWwU0a9KKJqwliLgaQQ0/7xAI+ls4
RvVLSREKPfct7DukoAw7GR9dT7Cg7bLB6ESV4Hc2KDe8bHQzgu5zAMKAXTbqRXQDYyvaXWZ5rXZ9
TzkFVuYeMAvj8BkK0e78MThJeS/iUNUK24ddf/w4B8USlVyGKCSiE0Ix9TGJzyNtTzZUaKJv4iDt
NEGsLFwlauXlnaJfuHU6A2FGI0gxwDtf7/ueLfS9NjE8Cj6cQK72lxoIJXrqVUpBMm6Ut6B3klwl
4KuIOKID0KkBSgCIgfiRfQu7vZJf6WGFntw6Ugwj1PceKq3QQ9NBmUEpaBwq+pPhRlMV6wlQ+TI3
5meDXXe1IqpXAObbQe1rkCaxPW3KsXiyMtIdtnx+cBzS7/CvaOkSRmm9XSAM/SG/6aDBWzvn8dXn
aFwmnJudpxJ6WqlOeFRVngwW3B2MKwTWNp6yOpIcIEoCwzyo1kl4p+PU2McoLu/2hzEVmGwOTABD
IS+puxvorxqFMA91IEJD5DY+ovfUKHsMlJEuqe28bLju5lVJErwhZLT5jS6cmAUEKXWVoasGMwGl
C34cj5OWGbAEVR58ABEyBVGBCSsAb1CA0bNldiGRakjgpKiq7Zb5myJ9gvwcCtkHm3GJFePWjr6A
nHlYmQszSZ+JRMYqWm9bi3T2midd0ZT4wgweTh3rP8KkWZoP8RYTH8TKKBhPWzEEsC4Q1syzYM2/
JYJIdG7cMdeCFKoQTmWos6z2yiT/gPXVUqBNJ9BPPR1Y/WYULp7QRIOPoIoYwCKktREFmKsxaja8
Lc5b6V9YcjX29OcBFk3++N503wXljOejiyKiGXpnRsT4cnaCPEix+9ppMHH7f40xseXrv36hQPSE
NWyQkY0dWhSyDsqGcdaHmkgp/FsfMJFVkUk1IeJz1ocLCS8EJ6vw1sAyQAj/oPpE+FUK+c8cCRjq
x9l3OybEr6mTkeML9arhme8LnEa0wdAVZzt6G9TyJdCni8XAEjuApFo5RXB9Ijl6leQQfnaWmUDO
B3KFYZGH5aEqU8BQcDmXq5+AkcV7LFGxjInwsjelTOFqNVfUqmFkyaUedHIy4KlyXg5v9Yc+9W7p
41h/9J2Huwgvr0zmrEk53QkSn9mgMV8augWwUYidTbagrC5j6HsXYa8Q7bdYxZ8AORkeK9i1L+/t
tOBGEbYfLJ0qQQ+CFvQ43MvW3SAfCAlbZSuBh69UB5Y7LJDGMVzZY7p2TNzDcnq/N/UmOMlSZoSb
PW4lzMUfoHbuDGMewLxubO2U/3LwBPNKMhSdO7JeUzg7ydsRQlrvPkDTItQozNzUW/88F4Afg36l
lhf8LMAR0P0JSAxxkfiD70eRYV/hKgfbFyNundKAFAokeyUiIcdZB1W1wPYuRB82UVvybqaGyQzW
RiJRDxdfzf3YYB4MPc0c7lJUh1VFs4gmIZqk+TZlojtW8YQE12DXGb0wJYiWwwtTw+j1SklgMrNL
NbVtvOZtG/KRjiCKilAvhJVowkpnL4rzlSuNo1vGGokDhD3pl0aaIMIp3DT5/GzJ75SA+G/QHuGF
m20nKKf8R9Ra5TC1d5W1GwXSS1n5977ZOjzuaIlYTr4xC8jArl4IPWasWoN3ZqNtnX2HFvMh0V3l
HUC+u4SX5vXRILdCiCq+qoTa8J4Ihp7Va4JlnOycYhDg5vGDHMw4+2e2ZZQp1Splvl6vtMVhvlWR
FkQlIGsKiG0cRHMd/hYJ/fZy54IEvomvG5T/ELYP63BZyiTvsOQl5kZ9P9Cu/B7qhwrc9S6C4FmX
8xWoIw1z9NJ3hgNDw4V60JVZWP7jI68Kc0juDahuTOAoH3tCG4GaKl2OBVbp/624UHJEWbvMxdlf
HB7BEgYU+9+BkhuLvoT7KrM7zYTKfnFuo6H3FTo4IBIjoM/WjPXDAeCAuIYcHMFbfXxDvC5Zz2WI
tgooaaqQSn54JKOCV4lbkqbfx5CwDGIE0h35y73/NpJa+O4oiSv14TLb8UmXFIgfv/h9OHP2wa7m
reigcPw7kv3eBlMdrtsXxv5jg8EyxIwgOR0qKc1UZz8bY8q6lWcGTe9DsG/qM+i3F7XRFO2aJXOh
4FtaKcQHkgr2jy869eiAYfvT0KrxmqmndlvW1WR5EjAAfZ6t96F5RHJTlQ4/+PyWi86TBUSw9TE4
ml7O4gwOHtt6KDwjO9yFriMkfD/6J1p5Gx8LU9GJ0ZshdnQTma34UNeFvusgIXvqnrU2vcLnD09w
+bkDnutP3yLjKNEZj+KobS7z8uWj4U7uWs+rXBYICgRYLzEdZz06kgwuJxASQXNAAapt7gNtxKOk
gbo8ezIplr6wQA1HAfxBDMeqzn7juJc+9zI5GJKNG1sIb6tXEJzT4HiJaryOIocqhAxuF9AjsSMn
21JYWS5AWwgMmDK6Z22/U6nyaWVst0LO0I9ZyE6vxRB5LuppVfRdVY8a1XcBkSx8S8UcoCT84TMg
405ujAeEIPwHdlGe59V/6sACbSp+YBUgkCyBpWkDHiYtQ9NA4TCiOQiZN6O95Q1UxsLBQcCwLB0j
Qp4Y5II99n1AAOfeh4tq2eqSkemda7X5GEMbxcO0LS+IF43gypUpDp2G72A+3n/tqDgNWavdWiOj
Ll7oaaSlCZs/U2C2cE81WfIBiY1oopKZ1fQ+cw+re8bwY/XSk+n2w2N5mvz1keN8qs8DEsbz+biX
E20CFffz9IoB2eakq04d0XqYrdfpAuaJ9Su3nnG8fzXjz+avyZAui2yKbL1yHAx4MuighxAgNIXf
jvSbXZ3GiUjdx8ek2SzL7WZNGt+sJSyKIxwiL8ZHInw+0WAGuNkUjzQnsnoBAwffpqLrltt1Vhx0
wohTq9zHjruXuJubjRkc7F1S8PXSO8SxZfMuTPEVJHSCsKAv/In2EX8LyRGjr+YvGkpMPbiiSNKk
3XP9fLoxhgzY0p24hr9lTmuSY5OeT/fOFnrQN9XSLGEXiOaTo67AEkgl++0LQ2RpzUs4JhF6SZRg
/yu1XGXR/ATyCynessgx5RphPkg0WWvreVtRPk03bLNr1Cfjnu90Bn7F0nJer+/wvbEks2AioNEB
w2scx3nPizkMAqhc6sqBhdYVR2qGYMmbbAjdkd/2Kotf04KrpEYekGSZHTrY+BhkFJxgz6/I6Ay3
6+M8RLuQk3pouXFqov7OqNsq56x3+hDOtNjsVo2Ev8d6pdj8rKnOrOung4zyY5xUeqgwN1icc2wI
V/ueoAXD2BuiCvAwgFx6WXASwzJNlk39UFyXhRPRzDxVeB7+L53btmibN7kvjBgI6SuMVCKBa4nE
FoNkQOlYmH+4w6WZNEiT2qwtZYArAkLVFJG/byI0/aXzr9VzJulTII9ucL3iNIP/1TKgHnjnHixQ
d7A16AR1cKowCm7Fq1SXKT85c7IPMl6R4ai7Fsh00mKvG4V+aKMnGv27tYqcXaVYcJg7ViUHSDm2
Kgic4nI7zTFkoYDZLUAo0EM+0v3Izb5FAtqusFSBSO23NPPrRTLZD9j4VaUGg5DxtfqOM2SP48MI
7a+OBw4r3EZg1+Pl1lIZUhQsSwIV2bPmBtO6dH+Q+XySLxVYgEEr/AngQtQfTwmrXrPhZjYDP58m
gt/BI/D7gNjFf3nChP6Cm6fjGL/f+ekgkU+J06k+deRLRxaKQ8LynAis/jj1l02SSOifgLGcJJfL
Z9+munIuFzxZb47nWsbwiumZgz53BBxeTyjTJL7LT3vsYbiPRU1EBKnAnRxZuaNqp+KejyyMQ0RR
Gu4qkQFoPjC8xL0VvJfP20UGeL1IabBnPSOus0jdFYErBC6rV9J3RrujFBOq+Grqy9bG+chrxaFU
A8QfBVDrJhTaaGEo7EDzq31k4qPx1DZi79srGoiJXSYo6hijTuZDdDf0cbtYMtlXjuo2e1qRSr8e
bnEQDjSTl4OTtEb8nYgY74Ca66FTNzr9ypckPpxHBV0bv4Y2accd85TT0QgU5g3NpxIBwWccJ3lm
fHzFYpHdg/n471Mt2tALsoduTDkP4aPfzlAvyGDf3fKClMDGU0Iqca/pcdvsAri+6nzqVdEJyH3a
zyT4276h2LoxBVMR6Gn6Y3oPkIlZQCcSuoJp6mL492SzqUlE6UWJPvvj5NrRifB02To8LBJ8EYmL
JDC2zCiWxosJTS4xBhsfDoYxNJf7/iFOR6zTlJnEAU8HczkqFl/4bSGWATPW4bSC93yAiMUUijTn
WzzEqqR9SJVnWTw7H15bi7qNllF/ag2zCxhK4dyKzdmpu/F2KvbpYp4VseaCNihXOJOvp20bztxw
C7fClIkpZoROt2vL+hmxCGPwHJPEx6viXpZkO4XoT8fek1WDYnylA2FvqnO2oJ3imRbwdz5lPTEE
tSZ76fVdQRgf/HeuMfNdiVgXy6XdKKDmzmg5PvgHIA0TTwsQ+9tHPv2HwuTDVo3We9y/j5rU5qof
t5MDUJP4uB3FkvV9NtNNV+vQY7VeusnbnHy4hFoKLrSNPbDtldGtmVr43ZrqKOe0oEsNEhDWgWIC
E3IpgkkBT9V6rNDkFmolQXg7XbM4qBghOAEDHuZhEBZrXuj67k/TRTWh8JzHiI2Ew6L56hfEUQMC
xR/L3QoZpdYK4mph2x6ObI8HnYynL/xtKOvt9ZOt5+SBy2zV7qlvcx0SLgM0mGzuOGe3/nSUvfFQ
EKKQqB/tTmcei0MIhesNHNnfCDoPNLD3/X/96uG2PAqZ1fBta7V8Q2KNW7s19lIkMQT4+44UTVo+
xBJx4sgXb7aK0oJwkd6oRp8l8HmhjeHFSUHVdGQcryiDMrxBV5cv/nQpflHj0imw3h9iGjdfBShF
12nmKzEV+PwMryFIqxvg3eFRdL99Xwh3Ecqb7uqnw2nvCOecjDVGZM0DXp04qAcSk4lQ4ZQ7zyDu
IAOSxB5PY2PJFaOo9/+FzQtKwWLfIZFDg6he3cYt1C0n+eRagnzQ+21imhMeUMz29TnZ8NkfyN6x
sahjIb71ohpaIfR7oWFVBlZXoIH4Oq8HsxFXI073v3falFUvUCspOP1+WSwXf8+huEhtgCnLgZkb
NJUe+1782GVyruorzjjLr+5d8kbovQLNIeHlfND4KPLAJRdM0OeEpDfeqACe9Ib0AEMzc1cK41Az
7IyPxczPxfuEfqMrsmKZqaC3WOeYxyhplfhzTy/oDjY+qxaKbjbyHFp6Eo1ENNfhrKnfCZIUVd8I
uDym0mXhzAe/1FenIgOxnRoTn9CBJKYADYp/BTVbFOSPs1tjsolD7Fx9GQUaKvtP1G248FdP9YMp
w3T7hjZ7rRMUpU4PQcaT6R/stp/CrWlQ9b3azlRkpbV3aXXkXCChzPeFowPlHxzxkvPNRRZrRJVA
49FF8nB2WCved6WKBRU012j4jTfuGiOMJH7YPqhNRy6Qa3e6O52XeegmuWPBgz6fOM49yVRZyDho
XsFcHJER65N5s9jtX/LducZI4vxWVg4AmJngSBhXkiQ07rMyZk5/AQUQq1/B/zT35MfBFYGUD2ER
IQgz0L7KSBycCl8iC8uLOZCiHEfUEQRWzyTS6qfZECEaEoS2nmmdTaPGOq9wKdACajbsh95Xj5MS
nHGM3nxmKWyy34qvzwAxlN2Bm5bRoxkONTXf8rjc5GLspyhdMZwrIm7ZCgSc0H6i4tvjNP5vPOgV
Uj2ri3FdjoXuZ+yw5tbBBwuMkuplGAr5nPuENsBVI9CBqal+nGL3ytK4jOs36u7TSwQOqljcXmXb
IPXZuue6ce56Oizr07PpH4XzdX18wjNW+tUSdoWlEQMUMvOb83Vv24IfSCoa1Xf3ySTRxr2RPDw6
Cm1pfwNPHpeJz/r78QiIorcIknWOvrmOWZP3Gt5OC1kzBM7nGGs8WGCjk/Tvz64Id6mks0Tn0VTE
3FTlofprVVwF0TZqDvR6TzoSATnW43HJySIGnVRgmbVleV7CIC2XZvEdogSF8v4QyVqOC4USsW/O
HcN21iQKG4mEckmBUyNr/FmFjIiId4iWgjMAyjbp/kllbCwGvCZSKnlAoV//aRa0YS2N21M2nWx4
C4jKezO4o7WluvEZ54f8aDAxcTFQKII7mBsoW1kRjrUy0OmT5l3ooC8spcQi7B28uuX9gHWp/Xx6
LRjyvRns9fNEfKSdOJdRMyxsODrhWyvNwcg9dZRzUfkocsdzpL8nJbTvjYxW1ZuTGOIvo5ZYnRNX
3i0hy95BpOytJZ9kCRYGciV7wHEH6r8w7rqiZDjBGRTCgreCmVn14QqXwnpL3x6DgRMIpKRYecdS
dGkp23+zmWo6Kwszkk0goycq/g5UU5zSBPYcBij0bPCAU0d/YjgLLA7gwOODWp9/Kz/cUrr/IlKP
1UmqdW2oRcQIwI5Hh84T3wVio8DPGsmRLaSu7F64XC6+1c7vU1XJzbA1dYoZ0NF8c7/pbpgQ597t
tX65jGZVnt0hen+FWi5RB1G/f3DyYfp1LAFVHMjpHIEXQnWM/EUKtTd1XoXE/HpDxAE9ow+TBfzG
Eiw3KfXnDm3mGOUbTO6+jX/qTnhvvPvwsdMzFvKoYLaZeipbJXy2oi5xz5nnQEUhuxmASfPg0DjR
rHcZEX3yBcUr79WFDsMCKttP0RzznwA2xkBA5wPSW+r7LEvGyxQm+5kTao0H+BY2jNR3qepQsQeN
xIPsVzZI64n+PE3zkzkbDnVhm6AcEFqa4k6hYCouPSbwtdB8VWjNWnGScgHDVDQAjglbgqWk0a5z
6mSTBv9u4rLwENrrk7e1otN2yyZzZ6zw0j+8/yqWoWBrSqX7NZI5a0nx7fooFs7wVWCDvm+/MW70
KrCVWA1lyku+iUId83S9JkrDfLCMfzaB2IqAxTkx5HJevpqH1MfZIi88JcdCv2NY/1W444piwN8H
zHI5iA3biEJUZDPlQyINZJ7slrTSKPv/LJxdbPyaPhM4k6QhsYAWpuFaTNXxCCEddbH13wR11Zia
CBpwHFSTALcjOr/OBUZgOyvrd4OMXX/id6JaNlVl7CQZm6XmNHMs144EMzB2Kzun/pB7BQk9Lo5j
HX9HzWrx2aE6atT74D9i87+aUh4hzXC6C0qZYX2u2PPU1yEF2BKLTwo1Cytsg8J5gFB9PMwFhGW9
myFp6uNHvzRe6bY8DCgARQ+YieRPnOwC1h6HmkY9DqMDBrDopfPdeRsDkk6OHHfAdzCeQyfbpHiK
6tI6AtU5p+l2HUuDhO3GVWjApyYg/Kq9qX0S9MLUy6TdgAgY1Tc6zlt4ji1XITXVp05tNtiaMUlA
uPNgiVPCH+WWC52+zd80FFzB21NKkfJXZ9qKGUeBZxzBnM6ie9D8yDFa5vKLl3VXJptCSDpM1O9k
GGjz5cOqO1J9+KQLFYyRClCN8vx2jckuDfLbFyjRg7oUUktz6ad2U68BrWSgxGxN7LUpZFMTeK18
n76PnAtkOBaa5In4+kA6lEQvXckYjfwcgOA1uNC74n+fHFIllweK64j/V+8LeP/fkrM8eeyuCFXS
TdTOeUWvb5o2OMWya4aX8PW6LdWV3ygSFWuu42mMHupA/5haMPv5DLeuwA/ikBL4Tewg988rWwtR
w/WOsb+a54o32R8Vj72LZXAq+g+lqIGMQb3GHuSQiizaRB7pqxp6YEHTZXzmxoN3ir3DFOkBuh6e
TNCK5r91wcJBRdWovTj63p+Gn44X/f0jkR4stFK7ZAsd3cKvGpGwyFeHVo+bkJR++VtAmt9a7T2h
RRvKNzuL67gb3IBDgb//LTy4D/CqlQsxVcZH3E0LIiCDajqVOWjq9Pt9b7uWaiawVNffkkjmSPgc
oiNenLAQ+gE/S8T02/VlG7VZb3qEXTSJIeqKTVjXG0ng/dOim6Qyjhw7otqkzBjgbuvNCAu4Y13K
kp27aLk6AKqGyd2SMwdbm7Nlf4Dsl7kvJ2v3Ktfg5gcnus+WA733zBHj8kCJ1HSxELxNkrxKbDuP
06CX5CbtSJM/r+58FsUmOI11ntWZtfE8Rzt6fn1OG16xawVPM4J85ORWu7P3OBqHj9pFbDWPGVGk
eZp8NuKqXHK9bUjonrcUMtkpQHr1s8Z5n8LQzrU6pSEtE9i2See2iEgTOYhbB8f1fl4bxbbZnumB
rKYepk9+KgIOS6RdfSg+iZO+r+p+k4T1A1FMA+nGgPSNYmBOT6vcg1aIuEQralPvu2Ozse2r00k9
AAVRZPHGkLQq7DguhHA0xtuEpevblTibG4bXvKRaI8n+vu+5+FIecBvxWSz1SbYhutx8bHtap7Ol
VnEhks2VxkMInel1Jpp/ZXsdus7wHB+B/zThhVaaAQZl9Y252MKoU4KBph5Hf5Pv8DsTyxdWaafa
0ub2Y3CmPx1JmJfhW7/Wxa8LFdHjc4WQE8jjLcLsbACBWdeTTXpS5P/IrL5DxurVyXNTh6KlrO2P
ukcxU7yvubHE0Y3/pvhE4738YL42glNJCykbVFwVaOfKW0GcdNDYd9BCaF9wjQEFSi7sSAHg7tfy
EjlACu8fiXgTNv1h7Lp+6/nBgCpxdm1q3jNkynwZbEUxGJnj79Cwxk6P0/P3MITJl5xJwogPiQ6f
grFKZeVXSibrCm7vDgUVpBljgzVOpWCOG/lPEpL/92qfV+PC9WApQLxiEDuxeayQGbv6l2KAT5Lm
60a3SKZLb+5BxD+jXc69dAMlz4PYtgYYbq2uetP/ShPNkoNgtPRpTzPHrbbmxEmqYqlrO8RbhAWh
K5ntnR6VjWb/Ct0aUXIjjcmm5p+lL4E1RJ1qPV7xI36RXx88zaRSr3LMDP+Unid3BB8W97kQWKtm
uGRBjuZ8peI4Bh1ML4+TLMX6y0y1PYnt2Q/Yp3a7ljSs+CLLg+t3gAx1+HqNZFVKW1dsufdx/bxi
jvq7DxTWQj76CqjkYsowor+dSQeXkOTFojmfDZagf+H98+0AJxRVBWN/GCptgkQmN9/mQBgC5qzf
mMn/QswE0RNI7dZHHcSVbYNWf12VqglrGGcUPcTns7Y10wv8vXBofLK/XU9RXIJn3DjqXlgukexG
/aJOIilWR1odar3d81h5d5zFotCD8jht1weWZQiB0VRE8qSdPqnugZl0qLs2lBPjU423CREPV9uH
fqW94Y/mLJ5yiB0AB5UEGd1vIXxdVEyDPDHpQwCPm1j9u/O+Gjzbct8KtDoO3mxXwPICWR/bPIWB
zGKqxc1Er3U5Ov4PUyQd41gUwqL0FVJMoW9dXJ3de4PoIEXu0MQg/N4mLRaD86Ci/O/CNOGZld1O
9NVO2LT1IImXTSvhAn0r/JqCQaM5t318es5FW50PNJ8tt3A+c8xw9rDuPlZgIyWXcuee+dUdrwwc
eEmlSNAulrxp4r93gVXIIgrgJD8uvwIYshXtcgRaSgMQfiLQY62OoEz52jJbzsoyPekapCv7mbSY
AKZ7qZmmuBd27Qxqys58D1gu8RiU8Fqc3ADBVLQkthv/iiAURDa2ifs6CSdj3p0R4CIOP0i1NIYP
WX5+s95vFRM7892YbF6S42m+Ekzmld+iSiL0gcz/pfNKSZhCj1hmnf16DX14K+jNwa3TTJUAOFvJ
K21qk3Q4/27xlYdpqKYeDaMCVxbLuRqnVhN9tCBAYd74jVuGrlRPZ1LCS3McdOCvyBohy84lrn3A
5qNDEOx/1LiNzFj5XInVZYsF/v3y2xtM7K0d29KNXLu2nR8E2aO91krh8DcKos83qLDyqY3Y0e+l
P/z+fgbmpnVpFzninpPtzoBnHb7GVGBSLWmNgj+X+vWCXSAINAiTnM1Q0MuBHjclRTanIC4zA5IY
uAx9JaVQ6sO5L6K/I/sZnqgu4ttlmeQNGqYsZgn7mYdLdkyKKvpQVZp1IEjq6mc+A24+RbacBszR
rvIRmLnMgRyE74hJEkHFtjkBfB23taXOuBDPg90K97EFhiTccJ3TC0SZ0BDGw5+LDch5bCjQuHMa
vjDFj+aWEIzT3mIJDDXNZiDJDOb4LmLl2Co+QOsyIw6fHFS+RDNWhdvaPjHcM3cXgRs07qA/i1Yr
LrNbEL+oiKaiAS6wydQY/zdhNJ8ZfbOA5HRgiA7SfVTCoPXP1Fk3PhL+grxbWswHO+UQO1Qim9tp
TMQ7yr+8BaBYKl1FfS/EMQyY2mxkOIk+ePhSb2BnkkIO0lYRDSO/5h3mgGTcNQb5b1/8YXqImuHQ
IrQmQdjIJaGDDkHeNcTuBGOKH+CsRf7BBmrbevx/yY/LeP88016j0tdPsLlObK5dKtydkMzxEK92
l3GbQ7V0IQQclmMWOEvYjH5EFY3Bqpr3Y3DWVXMIkFPd3tvgxr9pkIjWddY/S7ZiBJVN0rW8F/XH
FAhNB7sXfyI2HUOZdyPGysb+Z6lgOweTCglUyh6Z/1Zpk5EXWW2S4QT3RaXIszRXzA+NnbxR1i3R
3+ozkDyHgfZwJtIisQHVZIyHi9VLxnVs3l9vt6DsczcEC2+1qkTtG+bqvJeF15uIbGGRfdqMZdmc
7PNSOXrsq+eAHK3hGsbGQboeUp69MWUFX81V9gpDq+yxoP5/QagBFXdXdmZ0eiJKClaLjQNYaTe7
GTTj8t8l8GT5uxAGqBEUzFG5zD5YR4KY6uT8EMN49ATer02IfRvVp2PBdjI+vcEF7EGo+66p/T2d
eFAQOPFvyKkabqKyfK9zoP6cYeCPzJPEo29KUcSiUqby12K6IEl0/NzD85/LaDOB12CkFNYw+qmi
rnI5x2A/JwdQyF9bZuv/BNTR8BwV/4fltsTHRLjISt+0xQ7AgP3HPySRtxyM13kttHFBux7HtIP7
v/U1hgoGyFU5B7tP3e55l8eg81CYq1MP3NOM79tXeUuEJgX3QHZid54cyH11F/qlyJxlNxHwyJrz
xt6t0zw7flj5i1sHGtjTUJU4PqHVzw1OgP9eHzIezx/tDBn1DgXeJqeNnHbw3+mrNf2LpjxxibzB
c0yuVxzV3ZZy3MBAwhK6z/aqM/BZ3uZx47KeQK4yTpHVvusBFVdP0d1eusTFSuCU671Px1frlCD1
QEJgJGRZGpi+06KNUODahPHL0V95/rlEENchUsk4mBp3KKHIL/2VFCLilT+PcExSGePE0vf0nkaS
OJp2gVtJg729o8iaxN0aYbxASkg0FviKYLq+AlQnhNhDLmcscV9IFjRRhXdD2h9DVB8ovXm+ywDC
VZMy8FcjuPTiodbl8zOVnPxahPBK6iSLE5LCu5xDjJNHkWwrv9Bb3z2Ki+Cm2PhpOQCLm/A0oDrU
HqAwbqjdR6sfvXFeun2F0ujFdOFvmSnLeJ8YqjUWFl7iAyPewF2dbzDiHFFOV9/tY6NsSOXwqD6u
5j6Q/wTWk/Zf3e8PN+VU5iIrSkl/AcHh3VDFaYFcdOuBn1s4DiFon6OPu0odaPsXlfuOfz583ksL
syAfVIwrz8beZGoFa4ZSUqMms1ep9ZYg/uODFLLF9NIR/vJ9eluv3CFB3GlSZNUCtvXUGSppY9ke
bML3iBIQzJSvn18pXknOBybrWymSxdiw0rW/bYARV9SM+2reyKAHEjk7lZ1dUlZhEYEJh0uGnB9t
aO/RluSEMg9l3vINwT5j/LYz95GWQUywxJe4Y71lmpWqk+uwNbEuNhLCuXb+98TvohwbdFyOabSv
7i9zLzOnaJJyUh77pYjaN9vx355zckYHoecSH1Vq53pzfFJpUCo35kmefDx/gWmEkxaa37UvC/vx
ji8mukSsCKe8zVk9Um5HU+zdhuDP5U7xNY41Ajcv/oWTxtpTFjmrOr3h6fUmDW2FbgSW+8CeKfRE
sd1fJcTqGY13EmuLiBDetrQxjHR7+ztisYtUTBIAJP85X5v7uQcBg5BDTkN8OP8Jr45AV5NEYWKn
hVCgEO7CKqyqIa89ncZVM5Psv7M+Sn1OO07RaM5Z3mNx0YjTHmE1DWudNckH+2Ula17o1l3/xDLC
DMiS8RCl2q6c+qfue6+AbwattKQJiiZjwetyLRBskblzrwFnBnaUMmcMiJVGvyoNaAn2Mki14x9w
fRlUwyahhDCGLLh4nwQjXO7SiIFSlydlawkr7uQXn0zN4yq8Jz4DheUa5pBdszcj2r11wWmcTUCE
rQOj+e9nr8zLCE//QMCWfdWacbR/JxAzWSl8CpYoU+6YB0DmqE3RJrSqLo9ax+I5SnJmJEKMKQtZ
Z9k/I2UwncSaElZ/Bg6hDEG/UFccVq7qtkT1yH0HkcBQT5YV2H4y6009QXCs9MT3Tg50hgq7XNW9
fKer9SCZMzyCs9f7HgoHCtjJNVPnBsXr4r7jmTTrLIWExb/aRm4GaSdy5xP625n7oPn47jSsjamr
OPk+NPMg7fMonmk7nghx3725yE5+om5tf7F8JorFdNUDAg+7ZzFSzfiYxdL4Ulj3uwRSh600Sz27
jhId4/3QGEnterLG9NvKZFQIMYaEnRV+YEIHoB5OrEm1ORD7P7vW8oi4Q5nSlLFSyY1ClzrFZvbC
wxYgWtHwJiRfrm5Hoh1XrTcvYprLtD1XPdckXJ566t5nyFPhwkDkBhqYDfk+4wlWnUmiGvyotLyK
Bri6QRxsgk+Rj5tl6u89evte6gc8hQGS5jG0tI3JBw0Tf7fSUo9vibTUvDuculqOBRWl6tNw77Ui
qoEergin82J0gfL+naXxaKE9iq0h/At0FtmiL+7ugXhXdUgWWGhNmkJFxd2ca4k1BZOmDmbWAw8o
hPRwM1ZqmlLWNIN+XT/5ei5ehiENenyjFn5yCkErdVCX0qZsznq2ixAa9nGS9UqrnN7rygtkms9v
n6ZgxL3kVyXyKL9GIxJjQLmYbaX0SKx7Kvu3DLmX/4E/pnf9xtrOCUujQvJtZyam4BzY11vZ7jxF
5Yce+cixpPrK2TXR+77TwliKX/9ak/c0hBg6pNiKLGaGnkgnIZh9o3+5xr8+PfFH5V0ts66eEa33
Y+nvlr9VX6fOfQqdP4+ZKrX91la2K994dIwNFd6ioRpo2ar29DK0C2Xu3PgKSj8hR0RClJqvRiT3
6Mb+GL8VQN7sLS9CddqQZ1MraRarMiH2Ccc89LVDBTtOXZcnoBZzGd5zbO9BUDMfwT9Trr1ZeOHQ
UuH+dy5226ujzhfpAAl0l76zARJVqIasCjipZZ/EBXN+KzXykS5qNiWcT9OaWkxf8RBe1umm3rDZ
GDDnOCmbQsNngR3P9JtBvECKTDK62mZW2oT/lgowHzqwUrh5AbDDLr0y8an+lcAAwdwp694+NGqw
6N4IBIAorsbWmGzIQuBDJQ5vYStwjuDFRqj9m+3QjqUwd8dTnVEJsbwHDoS2rDlHI8kJLcyICmx7
UTmK8fuB/YqGcnvlgXyRySuGOurAklLfI6wFaBaWyw1E9Z6ebnniJ/fZciSONMCGi+HruvF/lx98
NxhrUJ2OJeGCNoR9n0eMat2WSQKBHI5Te3yopSRuwDJscHaes/NOMS70w6ZkJmBqKgTow81EvWjP
z5JDWjPdlMTr749F3lFdVpIe3yZhW4/rZ23pMqWWpLK7vgo7s+IIHwzaLNJNn4z+eoFah/7xX57j
lEMYOdeJ6DkYnaItJAJiR3DM+WL3MtRnK6REDZdbST5aC6H8gAAExU5gCMNnS5Ivf8PNyVoWGYv0
tLo0reUghsqP2lTcv75qNQiS+DFYq2IqTl/vNhC+8oQDSkiqhzN0L9A5G4XHxV4MzeYPmih0WxXV
npQ/YmGtn9hSWusQ+IgU11fdUraisAQXo4MPCBn7XQ2etxqdYW3QJRSChA4sHjY0yYa1kqDlyrUP
Nc9fvtg5wDtiJ2IC2+jEg680oKHBRwETJKp1YtNJ2r3Eub+VJzT9t05ldVz96FOq8ZX07G3vAIPy
Sacwy6Cmke7GRjmdgnFLUl9rE2Vrz9sJYkITy5EOi0g7TXUTX9iW2HcOIgYpUlbjcNz5RvTWVN0H
29ZjxmnIiOWlLCXIAg9WYtAWOPfx4Cq8JGE83P8ZbWGZgDXHXcd5RqliUGutYaQ8Kk2r8UiYcdjF
dBmAKVnVBbH+Yxh9WbbO73hFx0DlKUGGnbCCQf5+e9dCUxbmXy8BFiuyxni8jcIR9EfeyDm6GsNd
ChU+7vX5E4Hykdye7HH3S27gYPEPVeatoUbYjegwbncB1KePxW6CWfZlWcmhAwrSigkR0OQtPWac
sguTaBNG7rtuBLYQ7FabWpH09KWIkOy4yeMxBgwRgLk1FAoG4f6oBdX3B4diqOKkMEcTE7U9hqrK
o/Zdd67U+pzA8YkDamjHTvvkLjFbsUJZPKcrp79/8l/Gr+QR3nTJUkkZ11vwtiGI3J7uw5Fbp71R
WpqTDnzy7inWQf7OUsWy1Ecf/NpWoGaLF1v+AEJhL3U9PElHL9WyomFJD990NAGvmLcdP4kQywF5
gfTn60NeaaUWR+hYzRWJcuKvW28Qjs8gAUlrOTot9ij+LQB4ltHLtAv8fQzTTRZifTOnfaDsvRni
Q33K76MgXLZMWNEGOFgVqj1VvFfV4AXuNl34yDCQkUz6Z3JJ1gAa0DMTgRfNxpEIjd7tbWQ0oiFF
W36M0CrOTVi9RcgB2nnpfZsFOczTi+tJZbJyj4QhoEgj0RzGNyAc1IXSNvRrtHfBWlsrcrcqUL/r
WLRpaawTAScegyCCp0epgm0VcrgXldlWg446Qr2yyNsyfdwUpCLUODtqm/kIzP93q/evOIRBmcbs
rTI2O12ETGSOz2VDiyBhLeQtG1yorAdAmFmDdzFHpSwrqHC5iEZy7Oa3qYZkjIVped7T3iF6Ki3z
165ja4RmyAa1ex2+7+BGGgLYmMIGEEiksrBDHItFP/cixv49ClQX2LUU1EYvb1FP1iE4jhiAccld
sqaOEmsEAAWy+zU7KTcmfzBQNb1tFoXFxzbD6y2gBDnPwSTymTrVITO5RvOh1PTJ3Q305JvHvKLc
EhxjKGsIFWz8YIs4Cq5fQNUo5dXk2sBCX5HBmqNS3B/FCDL4tbYJNmZCnsAWz6jblvbPQ21AOvMi
XMr2+qQ0SQxWXtYHYEk2Fy9elkG35G2sT1htId4HOsRkJr80moWxJcv8HYwD/XHkXNcW0JdnA0dx
l4Rp64flaADkVRsXRJRN64wgaVZH7SEKqqnjFNSM5HQ1oUVHq3CKmFB8QeT0Zbl8qUmUB9uQn/Bd
K73J1yS3Jr1z9hWpNrPHGIEVv+oH4tC0BoT6dOK0xqb4WzGst+4nCQvhir3ZVaskATzmP9f66mWM
TR/ZDjJz4rhuWU5MgtnS3mIATk7eVjbR4pBj+WXyclnGll9UUMHqiQGYtDhu5qfqvnQcpwQnWhoP
GyCRFYs7tYAnmoN8T5pA1UWoglF1kh2L+VpwgUTQEsp6GcKAlyxakwfllzmXkz/ZLhw92Y06aooK
XuGCgL45ODod5zgPx/xfzoGYbMVqNVz0jpWaIjNAjbswT4M9KvNvo9uVC+faBFsQkfirTXZiOHBL
eEtqQcaQ+CoE+UTLaTwISsZXmB5LAxk/0h7NWkilAB4A9/+oZaPlGGLbL586FZrrxwgdwAqLjAqT
V7bbEMjObe2BrPL4Tqmw0Hcm3NOsZb6S3su5l8uQ4XWoOBpaelA284JyJHlmbYzGu5bV6PAkY9Hj
n638ELPZyHyqmUUHd6QiCpEpaB9Jhbk3D/MBKLKygEpl/pJmtfBf1+K54C2+erGPHoWa3Fys4tXu
uoryc14PgiqenQ1wu5E8bnya9TwhLrlbZyOkRLv/Zqy84LFMj/TEElG+h9U5BgI5Cmc/fr6W3u9P
k14YULI9bL5GZeXOA+1oV9S8jJL9L1c+W5oq6cncEsjmyKS1NV2aT0uiranao3MvL3wKp2yhHwoq
hpc8DTfUsHjiGrraqs7jZ5aijMhmkxp3gogHtvZD5ZalwMaNl063J3YkrK0y4P8NEfsG5+Hxe2ev
niaymxZEcr9cZ8iEN867Lo/9b5jjl4EcCqhtpi0+zCG8+C2dhEMLDR4/+ngIYuZOdytLqIeHhQlX
6ibM+XW+2ghMUfXOWHZQhKNQCxJe7nFB1smpYOwJr3CwKbXKytseNulC0N9gi88ZxB0qKXV8AKi5
PenctWj6ogqi4KpxiK7q3dYA8BpoAvN8uv+IPef90qR10ifWVj96bUNw+4rr7X0q8J9jp5K7/IOk
u4MG8gEiepCGP9OkyVWWtWw/40hfjPKG6l3fl+YJlriyIFWe//a086TNhQBRPjqEjnIOb1v4QMMk
aE+gPv6agS+p513+FAffBfEtOb6DV7tE3dPbOvWV+ql8BDG2iI2kDkoJ5Q7j+LNb9WdnUY1OFPj0
O3RIlaacCLOCvWL2P3eP1eafYD/YO3M1+X0ePebkLvI390Rx6QUvEPanJk/Wixi8ytJvhqO4Xnzq
+Gg6TAAVF9NikRRM14MIgV+DIm9G3rAvVyoIdTADckM4CcNTbGoh0KpsFUFcmnE4Ewf7doSYESRH
Mc0XNdiOYdPkNO39aCf6AQruelWQQLF4duMwovqxD+O7JK9bIlZo++fj5xue/ehjPlO1HQKWIsSZ
4QH4h9hraS0/I9ldigZKuuGp2SuinsDPJ68A6BMLY4E5L+PqVvoq+9vTSaeHkJ3HiV9kLc2wy7P/
pgwp4FWlxNQr9ATcKuEI6QbSxEKZwweF8VpYwqpZ89xBxO6aM6Ih4JClUo1ANeXd6Gx7ZGidUzsC
fWuq9YvrLcT2EswOL93/zx1tLf2N03iEpbbX6sosJolGhO4IBrA5piPceITpaTXupG1apY2M9ogL
F9Uu+/7cPflPuUVrhrZchbDBhu1MI+t+NA2td2qcK1wDiLxdqsMYaBnBZF7N95wCiokrQvCKTRKj
1+jDeY6qeKqBlMLOPCfIaDyU19RGK6l8HfmK7j46OVT9enbONhKYxU+O9Ou3A8rIDp0IbTs1AIQd
ruUbrU2bvHq+Vx+lVRpaalfVxB+HMDNdrneKODkU2BlQvx8h2dF6knO3WgiYWlIAf6RVVy++H+6F
iX7QYIvmCHPIGVTqyzl3Whp/RNl15uXkUaynhHPOkEtSrSDmW8zsyUC2Ap0ORqtnKMmDymi5dKeW
6IDHdjLnv6UAPg1W1bri7d/bNcZihsh5Hs65AQTmdV5CszsSqNBk4H75giJEXiwGA4dO3h0JxxlB
XJmrmR/zDLxm4hwoEJw42Q5UhLQNlRPm5bUnIoaIFvNncHOydBupBLbhjIS2yWMKEUR7ibw84mXb
9rXyWqUlD8kfYYqqVyaxqZ4nWQMw0PFlarzpA8PUKuZPL2OACrgr6xq6GsNBW/fhz25uj3sOfmKa
wICnigTwaoPH02TDpT6207dp/CKOW05z6zCZQy2jFrIffqju6Uv/p/U+FefICIvUJpdij4JIw2cj
oIm5zzX8bcclCVZ+HRfqKHpC/lDaUVFLUPsoA/ZAfoflu9FELs2yQGa2FI2tZLFXYsIn4Q4p+KRu
ZQmos7gxkKDCnLMFiyueYEgN2C16YVAYU2JJCSFfJfMl44739+c5ysQI+dGGQVRLDYhduvUBmfMC
XBwTkOJs8ZLiryD7qrMcINopPD3DvLSGWdM2KmJ1iUzDpbKzhLO1J4ecdvy9nXCrCqu/1oWZYYpo
jpml0dnGUngWYb09uga0i3xwf2UHLVJ8tw63eNuvAtU+c9dDwnfS9nfuXweqrh7X5/asAA8ODhKt
qDvUZ5Uo+QYFZbRM+4xTEVz6f4ZMzygzUDF2KthnnzFRdPwfR97S8ycvpfT7SFUNsVT3M6k933Uh
zze0N/PQCurb8p4uxC+2yucivdjjk/zCCVJo37a5MiHXqaYXogK6ghpBLsve3sKyyKkB0cZYO4gH
7tUaVObJxvuT1OAR6+zjcHm/RBItbmLq7r1A2cLo5XmREgklhmNT/a1zDt1iGjhC+c93GoInE43Z
GpSCuV8S5w3CYoswBjkIFVTKk0zSVmVBPY5McLJM9hcDuL0DoUsxJgF5EiVoQtQaPaTgqSaPeCML
+qQRkfiPTfh3PbqGAZdNSyfzHiVHdibmnOvbkSRyCkhmJy266spv8YFrdjeYSQWRC16U0NWi2p64
9ktMTKZZJ0eC+pb3TBMyfdRWamWFsjqQJwoonnHFBLgP37JYa1/OZ9Cn5iSwjwiu1CxRT8u9b4Wm
Y1XyyWioK6Bq6YUQjYJEj51EyZAPLtLtArnCNimK7OvovIXYkb9DgVKg05Lgyjk0isFV/mEmAR3q
Hmkt6MFkawZ0dRqC3JrUE6qzE4LsMVstOFY1+uL7PeUlEhCc51+G9WRh8TU8z+y+fe9MeRjd6A1q
FBoXZ1+JdV4BFxg22rJm2Z0OBnOcZ+BaDlEoLmHmk4iIyrGag4O8DHUpDxk/ccFuGsLWmOYoYSev
oyjmc/c8WGVADjJjW43kXMD3cOYTs8gaY2BCEgQTAiQ4DunkRJ3TucQ8nh8RKdGO4/ioziapcSkq
WoX04t/q7p9IhQieC/o4AwfYKIwO6P6QhK/vkd7IapX76IxHxlBTeuOQt1faxJmNnlcYHM974rBE
wEWl9XwqvT+W2Ke6bMF6tqljb4yx7Q387xPMpOZCuSV9OTbUViPBVJAgzs8K56zAbdK+az8BoxSD
Bw3Owt58YKGkmkITBfFesqB4vRr1EePTAtQqHhWFxnDxG2Qospu4soYpYdxDQqDPWm6c0IcJe4eN
drOqFdk2k6RmialwXPEplMU3BnLkRj5dYhDiQXZYMtzjLItH8rwPVu7L8mZ0gwupxebiiNpcJpOj
B82zYtX/dncHlD5a9CPn7WOiOMk/Lg4Ce0pJ1PBfMkhyxWOEHIZ8Ec63DtymGATd20D+CnCn1cTg
NTbbU9XNMs/RVawn11dBC1bIKoV0jYV8xZIdSkVS8LRku8ROjrNBJxH9jvWWefba6l6i1JZyWA3f
9HxxQpPLQDBSYZ9TQsWfMkT+bGpDFgnWHHZYCM1w8i3wEjyUEFPXG3/pCjuvbMIuYbzsgh6Zbxdp
fIoFKqJX9RA3V6q+ztrm+ZCHibEERNEbYiJNZjDslaRv31652DrpqA7iSTYnK8NcSXCPgWR9B9mQ
Z3PsLgw66WkByKEfrt7+ymFrP3UNSPuQEFBQyaRWd1HrxWmmlqRtzIY4RhLGFGRCM6h9Pj5L9U+2
DGXzRvPc5Vzpl72UkgHTlJqMN7zb9+vW2lSwHrNvkp/i8aE6vpB3GJO5idZ+oj6UZhz4i4TTkdpd
xZJ/VUNjNYEtnj5dCLfL6+7INZ+x+GbDxvimDnoHp1ZB+kOLRmE8zsfzEWTNcupRfCqG/c96eb4q
p2VhZjWzulwA763mH1qkGlnjKQ/fBfA/WgdYipirqzp8ghF69R2Wp3NZMzk7g5rN6uXhISo0eas/
kuJ77METAl3cVNv1Lb9AGuZmrdNt8L8e5mJ1oQkR0KA/8xjyh4QjW6UlctMi7QWIfuE8qzBQPGXk
poQQVs9S9yCNt6jPAxWbT4G/JhtyJMP0CWDEYtrOUsKCOMmC3FK6VmDusCO3U5wiplKucq1KNcqM
XFxXsDy7xzrVKvMKzOniDi49KJlDqZn6cyXBqMyE8cAUp7tdL3o0Dp/4W6jR0SS8HDDZJppWWJM4
shIfKvKYwKWYKSJ5uCC9jFePfuTCGEz0LNWEJHhayU+s2fs6piRXs3hoToYycJSet4yOWKqxzSms
W6fm4deVM5dUt0Yil15IzIxb9WCBE0RRy2KJsbxCrW7JOrc0wAt8rwb6F9qMdIqTTJyBIR76KHVa
aCeyg+WrDaqRKCUdk7a4XhAwHShnpU7OKD1i2SXp91nQLaFJKgKGlRq3Hnu/ty39hl7qrvAvX7WP
dSPN02ffxAO9YoXKD9om4XDDHVqHXmWYobrPVXh/HPxQIOnIVLCA5ni2I5vrbi0D5nCqBHWy6Zch
HCPM2+rHr0QvGvB07Jh+MQ5lYdEeb8XAGIUvOQHrGCwERMW68FB537y1Va+dzYjPCkVcsZEXjn7Q
Xo/Kcww5Wf4a3TaXmkBS/UISWS5Sqx6nYmghiywUdcMfgli9YeWu0DatsIGLeKQQSQjZuHUQeAjS
KWwN476AlSsn1gFFCrRqNoNjLmRtVsztFQnhS3Ej5Ph/yIVpTGCCKZ07HwA2YJLp6XHTVoMJiV9q
culnriuyagx7xRN/VzlS3gWIdXiOCQbv6xmpf6uGkFVxczZd7qVTqrokQsKY9BfCL88C07tM7w/0
s023HELpzW4ImujGvLKwSAL9R1fUsC6Jj477aJ4CBF04/z5DUwCmbh703MfZJnl1Bz7iXj/tj5nz
xI7r2wlzcHBHyFcZdJ0joee8/FFIoS33muj45luFfL4FYUHf4JuiXu2Xso63rxtJhEUK9io8GbGX
PyVwFB+RK1WCnaHjrLTts5Q/GLwsF9tt789/Jj5XQNw3KG0OEtgxnDNJXEZGDjR2F7jPMVjsCmpF
Yu8kh91zC5vn0KqJ1lH4PGa1fitnFApDhshKK94da08N7+uAHHReqXLZCcCrtggGxuxoRKEWBUIg
xJ8diTbDRZhHaHK5FHqRQZ0YFyOS5ZbZkeiubkBMEZd/ARiJ1UQnWqRtvESyE4lynHkIcikJSlRf
foenUBj5UoAua7+48sLOShk480iUTBu/d7YviN9DkHfKgL+NOWEJpWbTOv8ECM5wtZ5rMkjxRyGn
+CVg+0mHvGl8wGN2EUr7D7gAOwbZYzm4RaWTCMbNpj7iNiam5WiNleGxEtnKKR8TanGBJcfrPVBr
jSu5SUsGlVumdcQ/t0miFE4ANmnjAldpph/o4WXI30GCpofD0UUXDQMOGMBOh49LVTOMLDWK1wNm
v2mUfR633+gqARWLMEW7PqWeit8Bhw27orAkevNwTQKfzVQLT+jqeHHgud7Z539fQwLw2GpvjHpC
QmJILAhc+FhGbFm3DhfF9jxnEi8wTo64Cl5Nejwy+UMyvDgm2QDS/WtgAiuyL8Ox6SUHuCOs0k/3
0N6XIbE4XFykF1YWuNrEgPNf/VIdsFYukrpJcrDPAQWcgOAZVjPoas1XIewDK1KggxFCc9q5IShg
VhbTYS1nMjGX645fhbRQysmz5m5ffi7KSBgONGPMd6Lqu8WQ5zp9H6lKS1/fU5SiMX4ZhczoXLs2
UZt36kEJajhPux6aTnHgMTKCkwQbnHTWwkH1ZxlR4p41unJa2FZzFSWXJKC3rhHYppvxzfoEXloq
oGeff16XfIvfjUhEqpKPwmWam55aFlbjYhKyJ/J/7Q5oU9xXGNW3q7FFHTT6XLfr/tlBmpO8DfrV
MeG6M/6YaNO5cbNTlTiNAoEa3tDCOvE8z3ncRmn5L5V1yDl1/ZTlnEKJC3bt2pFdoA4uiElxhETa
uEOBgbPNmn7V5leGh+SkYOKnKJuAd3wKwvsrW7i6OAdh9J6BvxDuWsdJ9q3dnnWkQbXmMR1L9W4k
sXb+K7OqNDPBeY6pJy1mByXzotlJbYJiRoePgel9XiaxyJxNtZ6kcQK5Ffi7xQ8+j9Zbx7zgCAlH
Aa12GmfLBKpdkzgY/+F5Z/4PRCBp+nNUr4T6TE0yOBJMb1tw/zbPh1jK9AnTV4ltuCUAgq7nafWU
6BLvvzwPsTRpKhb15ERr8PJxl685vJ2LAP6TzoueJXLrOl2+EzS1yVqwgmOtQuPo9PSAR4hIf/Lr
xJJmkmIzOTGKiuJttgGiw8cARSpOKwWr5Ndga7yBvBCDdYJzZXG0loJ+vlJjkAalXX2xQcWWPSWi
pSaKYvSJ14b31f+hE/VB4PQCSfOp/I6C0Rga0V8chXOO8XvaoHGHJjqS31S6Tur5dIBsQRrCC6ue
zW7KeWEAF0BYzDcscdC+CkFN0ShUnu737KXryV056xK9uGgZWhFOdldIcYkH9350HyZjBDC5/N08
1e2BcTv42f5lN2fG8Q0yIkXRkVm3wm4JpQAy8HxApu1JVYvgU6smO7e1DtLAc1Vaz/mdpEtUAhzG
BZeTziOba9EX8tHOrzgVlF8BjbQznWeUnuPA2ATAhf5G9KyRRK/wpQmxTsacBmICWfB1uJCmzn6a
UzJgGTp6DDxXrTURqrjahmLGDZnt+L7jKhkWmKufBr7/jYDKKP5PSlSZNDqsA1uJpl4BkkGRywsl
xUkq3H9C9sY4DUFxnPa9Y/yeZCtGKrNPq3zRo9UgC/mAufAL+s4IUs0UNG73Zqya4zN6PHMU9dVN
JJJNxwkF846ZPG2GiSFjKEF4ZfZO5/fLzH+7FjgSZ0yFUvgibjPm9iU9b/sPkbI/1RztDrv1BXQT
ALWgvqp/eDcoQrhUrerVzLq/pIoE/P2tq/6B56qcKhBzyLQcEyT7LoLkMo8cA/xEmw3D8BtE23uP
NPqKPT/8nNIf7HRQ4e4+dguBza3TxhKrEjUtgZFT3hrjMwFY2xq3sPBqfX71rwo36RE94Yk2IGv0
Do65hY587MRfqZ4ffkx3k5cBuKXQGCCuMo8YZ881vewiV9hZhHU4O11fA31ep1/3owy6UUO6/qRu
aZ8cj1S3FRoHGZ3pNuO5qyZIlv2MFGZFKyoJ7O4fm3ifVJZrp6BeNur/FFeLHhMsE/iiKSqRb8LZ
+rqf8OFXQm13YGa+zgNrSa3VJdYgIdUoICqIYl6BMuWD0UUmOeEc0NnLinPvs55fHgKL5ZZIann6
fB8+B6xCuPpPZ9vQOol+vNBaDKx/VskSpu75GL9IwIO9UqqxSCrQLQAi3g3ZUCTNy/pKc1kynQKQ
KkFOiR2A3NPOF344V+rPZJwZTKR0UdB8qenVoMAT9tpywJanJuQSWyyxAC6p2p+W2O1NHcNIzsF5
rNbEXU6ZRsIDR0SAw7nAHYQSlLPdiS3KAG7y9EB9PRgDA0aMgvfG3cK9HAfT/rzDSYJhTr1NmHnZ
FNa+1IQdk62BuDGE1aS5E5VVKOWWD5mxCLzxeKtM7VV0UCVCnOgQOjShVMq3bpl+73fEnPrs/Pnt
i8kZdtJDyPb0CFZJLi+3bs745VHgGzfCZVDYFwuR/zVUaKmDMabH9r90WZrQ8ZAeBZ+5tfaGGryP
8y6uYZdSuUoGH9ZDe/vO2yRiSa0y0qHAvxBGjdHWQa2hLpVLgxgVdnEZrxbeWJrsdts5sqd49imw
x/0nCBeWTd3E1YxZaPxb63arc2kkxUKXbwx6sosz9iGhzrdn6HMWjR8+/pKaPYvDbvlq7BMd9JNO
oyU2pcvVYM5iwmUrR4ssqID2aTZRVcm3D140e2b96SGZJ3Z6gY2yOPP3p/bpWir4YeOTcST4UfHZ
ucsTA5ShFeCAqMHYpSGX/4ZjIR72h2CJkMYflzlp90yiM/gNdCodq1cPATKF8IpXeJUCnm06ABNb
3sTP+8HUXexqhKPf/xH1zIYRJHVn5+K1JrgpeJLWg7cTpbftdsp2KyEnV2YGbnGzI07qBKipeOxy
uwI7I/wJL7aDxLtUbkGoymIh2PtC/OmF8BVJeCQCEedW8m7juXcjCz92zZQAJm9uIL3RWcW70D1P
citpy8G8iaHJsw/NKvBKinzFsgBf3VR/USZtMz9/4Lc4snevxd5WTz9oKRTJUuZ4a5WF75SSWviO
rImlDpQ+fa0xbGJA8dF68JZ/3ynSB4ryEyLk0J/8A1tfUKdTas1FJ6mdRRLNgX8bokNd27XpkXRv
Cza0gyyXzHjxO6eHO+LPYjRSNEBMV1YBwdS00njk6wFIJa0oK36xUIYPFgpYCCNNJUQv42ivk2Tr
YCExpsWJ4oSHjyHX4Ngeu7iccEJRZ6LEvxvPwuslpkSteK63EeadG5qgU+dioQTl7HZeDB98xhW0
EwETNTO4orGpstO6gSDl5F4JxRg5L/XuYLOKhoFDEHeRkKWWUBp/DZkIYt7AN6i4E77l6W6Lpcqg
KFNJj9wEfVea6e/H6y/pJKYpnWEjXzzhAZYey1G99JiaZp+gM2bKkQWrVWk0PANC1pBuJbsp6Rqj
Id9dIDohk0Mgi4PAbgk7oWjl+XB1JXmMQ2Mi75scjAakSgiPOySz0q6GDHW5bz/nWu4i+Qu2snvk
w4OYgyduTIRD8hnEsRuLCdRXcIYzNNDNuhNGNj8DkfUfFGiI39bey/hhRw7ec2/EjWd6vmApM/hM
/OSzAIFk9xvEThtgBH+FhOS56GoJoK503eVsn2Hj3B5QN4lpAw1k1Ah9ws+VULyoELh5dxObO7R2
mDfZGL7d49Jt98jgfToKRKvEh/wG0dE6PdYWcpWj5wO5TaZzAR+m6hNc0qvEWDUxbNrNo5LePdUO
RfidiiytTKcqffcU+fxEatyx0JWDrEX1atgRmPj2ie5fcRjjyDl9V0UZ3mEBdh4MN38ND9LF1O6m
wibDMfENCxoQolm5LyH+haGGS2brvA2Mdeu8xPuESrutB2T2XNtU9V+3NNycs298MxSeLHHs2Kxn
kvf5gaUSxLba2dA9hZeQWgbCDflkrZfEhgMhyGzTlF7LOW84Gb9XjnxZ0lcT/iV+dHkkhUtu/LlT
enkbVesJCp4x1smuaqtbnCb0ElwTk/9rwp1mwxIG8C6b90rXYuEwf3gmU8M+35GPix6+7iT9Zvsl
jxfnejlQJAq66bnvQ87q+Rmg1tLNMwMiLOrrMbvSWB3mbmOFKC1DImQ6VYSWdWaZw15P3io1bOc/
hUp2EtcCInkES4YxkrxEbNmAD9V0zRi65qaHXskd18sEVh/L2O80Qcyd6daDlFrSCMcfjckGX58b
Bh+vKwJqiN6AJMvM1wMeG8Gep1RY6BnX50q3YlcE5j9hEKF6gQrqxbvK1klXk4pz8xxK+6LakrZQ
RG1NgICGwh1YXO+usabH3HDHm6Ud/X+gPfrCNfK7qfeBE97yKah2iHpXWg8DScmOLWSVghpyNfjb
HAcLZngWsjOxdnkbSMaWlvwjksQ6fvldNlS+ByFR+tTLJPUd4tMTPT8rTy3XKHzpM0OAWl3d5UwA
OFtUZGtsXmz8OLeNqSIrhohSaTjxjfVHjyVuvRH2+vclc0ON4PY7X1+QpHgWxzOou1rWQqty9Eth
2S/7OVgxNTJG6TnPdoVDNuyqt598QhFF/YajqaOHVD4tE8ShmwIUtRE3wghbCGMQxjJRo/bTOXNd
BqLwr0xKOt8FJ7LLa36z5kwL6JWu4UlrJ+ckiR17CL6Isp7nQjMgjOlSIcOK6dq3aQXlpzVLvNNl
ZFILDa497dk2CvAxx0SKkmPi/HFJY3VICZ9nvn1w1YXUaImtb3WkvsFe06Zm9i6mgUsl0JkPm6G5
CXc5iOzVfxqYfepIBpoFRNEqk0QoFFYKRAzuwFyK/zPvcdVJTBOigTi02wAF+sG1VFIecBvpfqOm
cbq3X/PnLyQLinsf5LBv8rNNZnTQD48T1hq8/Ox1B2VTQaDV1qbpl8LM2gFOASw7VyhzfRp4mjs/
UGYwJW/v1MxvcCmGxlDXKDQM1ns/AWgVg61ZD2/3eSyBwnv5BjOIgO0hywhvCv1g4E5Eb/lWXlPM
T2KbwOJ8hqWq0WiUZUU86TvQbJ8klcr2dlv/XrrLyuQHXiBwqcj87/6wNn4Mnod0omcB4ps1jmrG
LUEcjpOgT9SGHaf4PU/9cT7nuP3S9xL8QIThU3UP1/t8ojHrXW3O+xHXJh0HeDM9OPUGHeBMl0FM
6WXUKa/NCP3PRVg1nmi9fVcG5CxbqTSlT7KRhTuqLSPI1rhVZQeFEHDdfyAbwoO8jel9L98CHOyo
0EuUYCFn7jPJ4Kh8xMEV0LLFH/YamPyraogY3ZHyUBb9BucXb5BKwI55LOk7pnodcXT4b3OMMCoY
sYSuh6GxsXu7CpiFc6ZWb6G4cjp9EBtmLG7CNGvfIpQa35WttRhL9TyVOhzpR3LhexUcppu/S+6E
kOSJjmhP1oCBI6tgCLrxnZWv2dYRUuSUwz67EMpUSQUDf2DPmCicqMh06Ue/sLrW4omP+biE+rg/
Vku168mIHGa0IgjRyBcxv4vc0/n5HhIh4w4D2P8JkC6E0kWFo5RMvObtkp9MnyxM5iWWA+pIrJMe
5+qF8S1hn322JpXkexIydWiWkurvZcSSHlkEP3O2FcI2ckaeKtnuRGrQR3d/wnafSzxO1qjqHqMU
HIds/BAaZzbCTP/tSoIwuTlblvX8P1loafScn3Q+6gWuoZMsrt05RwQT5wZJwedAeCT6IOtxElMn
mBR1F8H12O/SLkGWRqryjipCpAPTrjMlnUFNynlq+mazzuE+xHJM8C/caOtqnQzXUmEIlXge7a6+
1FBzBQE+co4RnzYuLR5BcjTgnDbVeyAHOVVMQ5DEDygBeNcmBahIq/W0NmYkaswp0Q+Z7WgLpg6Z
uLkh+HQ7/vCEpbZqQw/XzjxlB8yegBFMrzIbVARwPNp4O0JKLJbbo9eaZ1uB/7HsVskUodR2USip
JwjGU1nEmP9TMgZ6KWkadxBNkYWWDdfVOvVd7ByHToONIR4xgy5sNFvZqfKk77E6hg4orD2/5Nzd
Ehzm1IM1RbYIqFbZM7EOGvv48xsh4nbqn+PalgRAlXWc4vL8T1gFqCHLGbtWWJhUYa8oszd+3WoC
k52V5ahkLMC0tCDoSRM/uShmHCw1zz6GOyz7UnLzeIGrcbcgrYB5kFZbX7MKPsMfd8oVon0EdvHW
tSFlcA+l/7fZJceh+soaNeIkX61XS8ZxiWhi00azQfQpe5KqJ9rnKHBde3csF/mY5Vrs6WC6M12N
siStpTFPVGp10OTridUNQI1PTLhZYN5x8YTd1sdZdjEj7hLnKqLtJ7X8bkwfzxMGxWxO569H41ly
32qFkHJji4IfRyNULWOgscmyCji3P7IZHWxFOUKy6kEwz5IF8+IX/mdLBNN40npWn285Dn5p7JKC
IzbXqr53PO98ZLXiQ2p1HO9UtHFZMyyc4zNT9ME/ZI2sf0BvWsROla9Z+gwP9E+XFJb+J/II/VkO
2K9KbD0TU6WTKHsCRh2GdKpjWlUQlOOZwouV39Ycot0BFntbPymWFcDOFoFu/FwJxgTmVdh7AW2K
Wo6XgWhW4v/+GCmEWf56P1xDekzgee0Cdilz4vmkMUNMhf0AEzPsAMy2vQw0Qw//ix6cuujBL5RY
5VpFz5Cvg7qwg4uaG+K9LNyGMpQ8T2tAQeXU2PPGmV0tRAdvcMxyY2nMWSDVYbYuEj9qAtdlfpX9
wg4edlaTge6+JpqkQ3TUDDTTWplaAE61aQN7XTncjLiaZdYr8vYdsnvDPH0vKXoL8GzVrVxdIUVw
LvurDkygvNjWxk3jz98RKTYaehtFIohwaJ0ry+NpxBP9bnOSLGO7C3jUJAbnKDddlqx93qHt28Kd
L4FbNWGJ3NOm7G3OROcJQM6bKf7kFiqY4fUWT8pxIwXlzgMaWqn3hs68yaTS4A4/hdD+/mw6Bl2k
rc5mTSjgpoaI6xw9tbG1+Co0suDX2JRosb2oo6KKTJ/7m+LG9T6RKq/r0B6Ffgw/UNKXn8A7dw8a
8J8GO+ACk1nxBzsCqOSI1BfDrzTDqNIwjOakkNGsqNFyY/sjbvFynZ8UPt0PIWBOgZ/xHgYnupnB
AsjSXOjl2LIUdFyrtPTnf2VcoPBcwlP4BtcxRALC9Z1M0Go9sm/v4ZjpJbumgiDiLIKGljF2xjLG
ArTp8193R0YX+Xw5pZ1QpZAJrnjxvu0eIt0ytRW1mxaTvcqbkFtV8GJdzGQKIAQz2DRndniWBAwS
EO899k6TnaYbaIQh6iomu5UhUCJSffrwhdEfMQc3JW2oKB2YdT5I0C9t/AcEsEMBKiiWwAj9jtCl
Nnb50F/7ZJD8yvF91wF9VqroDBqHp7SG+W8q4Hw43wbj4+HVmsLtjiSnGvUXGbaLRQztljEuMMoM
IhCnaAXlfxOg6V8sf/Jn28my+eOdH0lybKBBv5qVDR4va8Ddx012zD3831feVIS2dQDNQ+QzT2j2
Tx75x8aHDB/ENnuC09p9SZO88yrlquQmf5PGLeY3BOYCUzIfxu9fYaC4du2s9Pp+Uqlqo9HcQTfh
aKIad9+7cJ7pUNjI5pjj71a/24ySAYIWj6WWrOiHENBIcACItZbke3SciSN4XT4VOwjt8adu5eHe
YP63CI9dd6Y10ZrXQ8bZJCkmX3/Q23WMKzhuDsuDUch/sUT8kBLitFrrKQnDgRz2aL975ngq3M63
17LTdGoCDdHiivogOe83ZW7QycjEBcl3AXMsn0znQ+9HJ0gKAYou6O3vYuJ58jugW12nEickqp23
oNQrDwYUC7jg0sxmbGxR+tgmxujnJLNuGTHoXIXJtt09ZwXOTJriDwws5V1kMSjcjlI1S1FacpRa
VxCxtqD/Xl21UMUA2vUXcFx9YLev0wpUWV3C8SE4J4S23tfAI391ANxdgH2P/RxDdReW/wI1y/Ys
BPKvUpHunMZpADQ9zVCvmcMMyknLD02vm6H5wEtSN6ktgb72fAw9mbITtEv8TnEnjW8yqDoSd80t
f3oINiWDhtgcl6gB2OA4mbdR9vqh5Gmaz8VxYyNRn6+xe4TBxkYg7bWudKHPoRA7XFi5pZH6AU8z
9S1ikgMDMdcd4hFOpVzwZIfDbWj0hDOy/Ywc32ySMTNIfBe3hUaVdPEtPIOnM/0LYjCGiu2nAleK
zg/IvLGLLYc3D1DEeBzv51eDJGyxAtzOtR1cgpp3wl+jwXXzEftAipPiC6vW4szzHXwvA8URd3P2
x6JHHZLaMroT8Zs62mn/2PYadG3X0CxgmCmcXtR8Mti6DVfjcD6alFWuMRj1eocu/P6oBjptbmH6
1UohMMnrlf78hLr+Xk2CjLCYrRAOxBd4k14FNfsfT2OFhvEpyr364GZqZA8ynlRdjUmPfxlPnahD
rF/CkjTL/t4dGCh/A+eZQlkat2aZGrH6FWYkMDAge7XU/uarIc1ZcBbWKovsRUDrsoq8OhJXvK3L
4IsSOWgfIxDPHl9PoHwTMFYziofkkMcf4yGvekiStCeOuzHpakQqOVWsWZKfFRtXbmLop5suppp1
FPZHy4Xs1/mp+9EdWgWSDCKbj1mP0Y8zJUTiiRCvmE1od3KftQMZKRceqFN730nzKvUHs8OQCin7
VQv7lZkoNIhkVdpI2OzyOolgl0z6Ldskvy6YxR8AFLFbzndhRPu9IuZ92gWVLZ2yq1UEH6n9tZsD
i+Hbz/6aM+GIuuEubXyagM+SEGBFjODPNuvmmCcxPm5LyZgwlcBAtlq96Rq5iLLTARTJlsx+3csG
LEonJN/5it/4nq8/RnaXmuhqAlzgWxQz9VMEN3/H5u3ikqgNOmsU/ev1dF07a7c2kgCJvtnESzQf
iFxvqrNp9/2VelJSjLTtlq0KdLfsh7nDWkFpaCSmxOnwbURbFnpn5AY23iL8ma9tH5ekOLQvjTOP
Vw1gWw/2ByKoSgidC9FxVFWGTwp9akl1t7dwnb1t84bCju1WgeUiyq90/LBW1M+xKciqWitIkN0e
9FFu6n5HTjOfONKcChXm6nW3R+6s4cBtCY0WI/37lIzrWjJCduPAqX1MKmV5XF78ywoK9dzQb0jF
C+eh2koz336J5pzn7AWz9p5F4Wqszyw1595j2F5o274iLkJUAOiqh4TUcZ2w8xnWteXLn6Edf4be
ffhdBDAL3rUAVD+3bJ2mzQ3v2BlIR1JP3yu6bO8r+Afizj04gLxhYyes78DAcxA64aSCpkkndg/j
15BuUwDkkatAZee068+ddHJfxPfECoBULkiD8WW5e4vnMEWPkNYZ0cyymn7cDaIC8rCX+HoFFMDX
I79huTPeVHPS3pmhE2xi7BnhJgx9+/MOst7cgPlnbdCNB013Ff/JywjZN3VcylDWFEhJtZyOP4+T
khpJrIPQzj0Gf8u3uvJBwvblorTzR+PjQ68Gpu4BCBdBgGBYoWS22g5QiAiE74xfzj16P3yqwo0R
ZUc37NFUAZ2MGjqYorhre1VBNm9egl1P/Pe+zpihp7H3rcO5d+uWmg99ImK/3D95GsI88NKnNd0M
z+5uqy9yql/v5d+/yTcvG35Ymvdu9/mTSIoLgovrUIl1LVI6F9Vwc9CvJO+9YuURVU7qAcz8nuxk
ahi3dGoqt1yGJ9CB1nJvLKrbnllOtmWoBr4nKZ6JVNx8zP3NOIHSeeHnFTe9tTmnTovcfwyNQ+Gi
q6wWqhtpUj9bUFHDgFf/o/YHaKB34Bcr48WHeihVfIc4ry6LEwwa4ToZZjgCjNmGN8WaPp6mVHa7
Zhmp7jYq2icr0GemGzUg0Cj2h0sE1619AlKAwDhgqdicRZ0k6mz0XySZjnXvN+vF6NLf7IS3vO93
Jsy2cAT9JdIjoTXwSN9axwGSbeaJCrJc5UiEaQCUzKBlbB4XN8Ppenscry7aHDJxGos2nHnGRyLf
VxoCQdVZ4NOikksNyrmvYXb6KMFgd45NcMhedhnRxppR7EWt1niQDgneqq1OgHfyu2EHUirrITpd
egvXW7FYSiM0dwQdmdGnoU/IH17DbCzarrNDFEB3n8s01bs+BVJNSJc6G3FQs9lYA5uHF1Xfdo5A
GqBmqMDvKuikLDvqJkUuH8NNi4Wjq7duZ58m53A22oLcZchCsqzY/HK+sSjnRB8OKt2iuox4qtis
6mNzRNh3y7Oz3SPGUBYjWgRlEinjRDl6eXyN52uO7ftwHoM8WKZlJRccqunUZBEIkaMFjCxaaeHE
19KiqYAy1a/RSgLnSq5lAuWtDeBZIZytz90hu/b4+fRD3ATkL+uN+LnXZeFHHomcUQHnjA+veG0G
jJdmEp7IhzYF02eDpzmD+XeS8mHmla2NY08qDESC2BniX/i5Oi2g1SX28kQFePlHA57CNjWxQpv5
yaJXUl9btW7nJroN976xZIR+BDMUTOiQxTxzVxcEZRaq/Gd3CHVzs2IWAkyfaLv5V3ssvsL+eYKk
oLFaqdzHT7HJnU+JarzbbH0Y1b0wcJDrun3ShRbFkG8kIqFo55Uw/EKn1Na5VnJyPy2u7F9qmG6h
1hEglH6q5LWE2Y4B58jDdAUMDb6kolin8ckOIuxL6i9BVdG00WO2PcVs7KCPAhs4MFadLmfdPreJ
IQ8d8shSfmE00xq5p8kz2ka7rbjLy+IhBLznbRaPhUphWZ4gdsUV8Y4ywc6cqMCYbi+jKOVmugi8
5Z0wDtEY5fsjDwpzrTgo5d1Nn1Lgc/w+Ig1HiYS6a5lfQ8biydvQqWoCVSP0Nl63FdkPd1BWzEV3
Eb6t1n1gx1lz215TQYmM0+cT/fR0TNOpwGWEEQXvl8cT3AOEoRPweHMJDJAVzC+lq6F0s0SFXtPS
M2pTIkqB6T73E6ztut0fYsHGwGp2tvDb6qXrNFA71PZGymoPVhomDwakTBSJHzTSD8X6gx+D5+71
9QsNxFTPiGhrBK2lq+6+IW+A408cELkp+lPII9+aWyNba1VmL5NTLVnARoWim//FhGHSVFlK9VI/
YXGcJn6zfUw0yIygxnaYXrNgo+ZwpXS1QNODQps9wWx/KJL8YlTegh826VAux0SZJLl9cIDm3EVd
I+OQgQsSTux7psNTofbFKCmO2nY2k1EhmX0WkAEz2GAFSUb227BZD793SBsskWN2Ls20p7Cw00iS
sLt+eEr/fKfNpcsXg2x84cFo5ecNgA6gZZUrTpNrjzOMKQu2hQo8D39G/SwABcSlmNdCzv0o++GA
PC620IpU4L6p5JnLxaVAWqB+WL+sccxVtbLwwxNKcrN8Ih9sM5EoJNCT8aT2KTfbJONnIFhQ5/g6
oEfeMp2yojKap6i+ilHoyHtUZqIUIt9iEnS9MZbBadyDEtZAl+fdAx3mi73GHFIFnIEFC1fIDFQT
g7MPkA7ihR6vQrd/imanECP8ZRdiUHjd6sqFOxz3A8nmeQfGxTOnIWLclfIYkOpUb6aA6XjwxYV/
Cnw49fZ53ZNz5Ml8y6ZxFsQ5+qXk6j+oAdPh68bKR4T8M6gwbZ/LE9D4APVZ+ZBtLoiF+9LTyIR+
kVeh4JZGJ2T/ohNvn4P/oUjojuvBHIfGY/2ZvvQH2y1KQSsGsdWjGb46bxglsHZPI6972C2Oct5I
gzYBrMGv4VXMZxH1aC9/maRMfXmbC0K2t1d3mOXhlwOv9kjoxxCJCsFvQBwGBBleuSM2lBbkWp0k
HCbXz7DUTrY76Qbjhfsrh12XA8trGWQtoR8G4nVBnUdlEUgul5Ifznr3kC1LBGP++Qx2IbQIWB5a
gna6CekiIAdtE68/5B7OsLtE+lO87WgmM89EVGj46mm/+dgJXSm7bfF+b7/rJ7xz8YlH/GQyWAMV
3eKm5MRCp9jAtrlqe/wuZ8nE4+WeGpyFlecafK+obEHeQS87Q0s6rFylJG3QqaNdqgs9xIl7ffUb
O0uvhkK8l3UcZlRvLjhykjeecryQ4fVrL5B56UzH1201/aSoVr5wghLPG9P6XyKzATv/rcuSeQcp
WnnO88mxQRutJJbWAQeEPu15iD/xkpF7brubevZeA5WpR17i7LXepWR5ducU2fsTBV/qC0XNywzb
H8TXhVA0HEoJfSaNBZb1nX2eE/vnppziK1RBHRZHc+c/0k+zu0VFbYtSzsWxtZwX4Dq7Q65KbfgQ
E5cc1UvTylZnJ8QDwvp6m3Kgf3XgT1Kt8Wkq8UyGIW7MsuM2ap9BeUJecp5Nd6Oy7N9w14O7mUzp
bt5BYFIcXZU5PE0zJ6ryiy8rr1orWBy7yg6F1Bu2JEyJcrBIUfkek6rK6KPNubyb16PcEgsHzu4a
14IlJ+64f39UqEL0EEp/95kBpT34jicN8mDmhv2qrkPtRioe6RRc2oLpt+eTfQYsZIhByEox+Nmo
CzQRH+u8OrAQK8Qh7kgGVmzuzYfyDpuo2SbpQE4GMUSCkh9uDK/A+HwbyaePp+NP6F3ZgAUMPEEQ
QadXW6o6wnsa1igwWAeV9q3qUNSNaOEisIExNNtMD7HjSdywGjBde4IKDwxDUEQ8jDRIHouA84dd
nxffCTm7XT4cq8hi8FSOir1YSBmMJ9iXT82Nhr1h/4P+AUutgy5IKeL66ujjwD0ae7Fz8HElanTb
/d6QYuYvRzeaXsnds4ouRdQ07hx4DkQTiNlQupybib7eMQUy9WudEMiunUjWqutcC2bqGE1XHqPr
Jy5xW1XDt9+rr0CVpVlCKcOGgl4q1EHolAqOp3NzLrNpWyZP+N84PyKQ2B0qf/H493mUYOnyH6I2
piVAzynu4u0lnDcF3YhqCIUXdel9RbkqvdxlXpuiT4WepM7EaWIhY4ix8ileOihHwOEaJSfe3trm
E6Bz3Q1AReEdA+LEOW2pA1WHTjBBqyRzDt7BIejdqvLl00KHUU0QQNDZHYQWjUFqjKjPYAXxOHUk
DuoUMIsNzZWwkpRtwFcr4kAaWxdsU/nB/QG+OM/0Nd6jHJ6vYhGVMd1SHRnPh6SrsK/viqK932Ub
o2MlE2pSOpTogYQ1VZDJguT4n2W7toNqm+7XuPrLZ7UvSjVezzrtRTMMOI6qAJPCzGtS/aDjPHTn
waHXHAbLT4A3TJ+Vgq1j4tjL5hi777jre0qVcYZjGUXvtz7OpPOEYZskzFT4q/zNul7gwzOXBnAJ
gNCzmEkpcnVC68+DKISuji0sTq4etmjgBKtWENAv7aF1KIv+zxbid9I0uzOfh8iM2PKLwSfz+jYy
PqYtGAmxtU08jRlG+tW2WVZ7ALmkPWRKXbKm8vcEDqauIUhK2gZVORy75Y09+8R7wZnrktj5pYtt
YCdNLmXeRbUmEL59KqD9JlDMkx+MjCjlQ37EKNotQ1EtEx/W5yg4l7li+Iv4W9LdGqjv2uj57cT+
jh/yKdp/mO/LnVyWJ7Tl9oCnI5hv+ymsyYcaZD+3n9uNUl1Loda/YR9jMu2Vuq/I6PKSZjE3hhr0
5opVsHN+DHKhUS9i2g4lLxRRjEL3YFhxH4w8RSf2fpc02dg6JNW6OLUFVN3JPaHfvmQA9+/ru+IP
SA2Nc7BmIXrjhBplUTmQclBfjA3bNRIow6FURVdKQqj9Hr5gvQM4dgB0iJLs/4G4RvSw0sy8eCXW
gcPcbNRAZcZbPEKJChjfOUtBTFzEL6NNkIkCXCF8ZT5gob0ceSR5NthlXQKr8zDKRjXKMnKf1w65
/o3WhcXeyKzwSSetH8uZMp2ZreungGnvC2JfAHJvSDdfANjRStWPxDuOGRHq8PWUjF7/X7gs/TRV
ewWihB7ObgjOpsMSBkzFq2p5YW6cku8XbRrldG0Rmrisb1vbbImeutuF702w2JC8iKLMTKegwDm+
TnJGhMU71Kuh8S6U7ujbKEvg/Uzu6vluqZlSvMUcBel8Pg4nrFpEBav+uFtVu4/aH174fYOHWkSg
O03Z+Ucbc9numtSeUXxobGCxOW0s/go+OkgN++KRY6Sl+4w/NP42U44625gIqZLxkcgjklrZCyO2
tpzka6QZ1q5KE74PpQhEJaW05/1hwg5Kugmh8VEHVghTc6LEFfqSYUVr946JmNkxB2QhHYHy7LkX
0ChDjEZD3uE+7GbpUpww8gNx6Lnu7hBZikE6GsNt7G43f860leqetfPapiOfZ9dNYqv/Hp6iJVlT
sHwN4VkHF3GQOmo3Ktk/kqFULclAf/C7kbsc7EL52I91DbeaPaifTQvJ6V0PrC6QKbTEtXRQAYEA
wVGCSnY5GiO7URg7+taqlmzBsKY6ni5fSX3taZYelaXOGdVe4I5RzN70WEuLAlDl7sYm3+jNs5Zq
afT9HAcBCiOyVnLvdgcaJNg8j8y9tBG57YrBjtwgpWrZ7Hxu43dhsg4WtSjtBeYS5Ppqk6h5ZnEG
y05wpJJ+bdX3kTxfq/2FF9MSn1xhta51ifk8OXkIcdYbEVhIlorb3w2ke5K4qxy3/D7hP0h/XSUD
s5LFN9UigbghHwAZY5y642QJr+0qjauwPgQkQ/3xJGGf2GR112zZwWvKfhhjIsi7NO+Jsh8Qezoi
XQ7uMI/xTOIxndNdO2tgMH7NoSVr29I8GzmTy8/Ghxa4GUaUEcrywqHKoTMu7LEZzaxJJzZZmqVI
A3TVA3TlKRIx6+EWp8h+38vVA2jnf+NyrCKk3UlJ3fD7h3onFnr2lDqVUkQLUk4OkvFb2eydkt4u
gj/BfziaKgN9N3QMIY0Cr4kKgzjdvYXFEzYJrlgrVWSnsqji3Ci9uYPR0XzpPv9gAybC5+3Eo3ha
B0pfEFlk+YnguBuIyzBJvv0aheE6J9x+xnXjaNRvFT9+sHkc9qo17GPnVf4uUJT7nTLjp/J9SkUE
ruXQb8+XGM/oTg4QHZ6OVNqc76pN1HD3tGTKwGCge8PaxrCd+/5J4++/VRiCix6tYi953FWoyihJ
UryvJzwQIU3CFOyKHvxELLuCddTYgrQ8qCdWolO/PtoQy4AbVgWXdXLd0DS+czN8QHtG7jDYz7eU
8bNwOu7wln1yyHvEZ1L5LvOkamDURJh7GJKwSUGUqS5YOs+tTh4xIJguX/rMufdOdjcc6OYbsRor
pcYYcAYKTXS00Fe8Z3PISObFvXtypblcp9SWUz0PYTOacxaSgTlzXj7Zl7fANVf8WJVpVVHOCoWQ
m7wnMqkS18vNpOmnVGC8d9lkqCONSeUm2CC8rBEimRGK3L+uDqXTuzyKCFrWxD8EVWqmihhXFMKQ
L47QPzk71ae3AsnIuaR/qciycz7eovIG6yzQZG8GksmKzzFZsmMwKQRpg7NEg1CrBasROsrSmpPs
zhfv3rV1CE/afb7+UE+BgQwUubV6gh8yBZJZ0vjganjCPBcSbPISg/NbaSfjQ95hkFkTGZOOdwt5
sb0399fP7L51zGGbCNKZ13PC9gk3uHLyzW/T4HekgMp3zWOtnPqQkGnwzqKaQeyyRwalHYHU3hvV
ozn0DZcJkI7LVqZD4C156Y6YUTCycDPFkCcyJO9vElXdrjVSTSWUYxJOecBAhg5KG0CY/H54SLsh
motcUNMt9J/hpgpRxLnh5zXUFw22yf/HSXXZ1p2NFGovFlSNnRvyMw2EVsQVrrrqg9C51gsNxiia
R8kpB6I0IJ+lVAoPqFHi+bY5c3hlRlHXtBDOhWYj17mFwlqN3yrTBwFKFMmO7Y+FZFJ185qvFnD0
947ATDuzuCJDhsYrVoT3hYgOwSzNOVZq0M0eXAgKi7kdZm9sTJGKFc970t/KpDCa4HkiVJX21reJ
Fp0QpMDti0s+fd+7UpYSIioBZDgXepgxT+C+1PNEPMZzhajqL2VAkHsFtlSV2ydMDjvB42NYhGAG
DFVh0d2qrCygSOEYcavC1CXYrvmDiQpKhxoHt6ImI4JNFCoBGkc/mh5slSScOJT4dBNYyTgoloEf
xC0CSiUjXHCVtSohtHKFUgraIYA99u52RSMb214hveRZVUTulobDuQViwlSKtVb0v4WkA5kpXZSz
rXDaH2cp/NBOL5pq3eXQnyAbqj4jrQDvQX7XT7Ts2q+32YsffgUIHAJHrUDLAR6fkAtWtAuraPOW
aOPgUeV31BOEbH8DtYCZcu7J6oi7aepIthkAYEup50EGYTVHcAg4rFdfdEIx3HxMKabKEWBAYqFv
3oHE5DuVgoUdDcXsW/o2kBRNhE7h1iyqPELWBMzwNqGbeoxcKGJV7MYZ4fHLs/HeQT2c7VhMJrl6
vzBnBeP4KM+MQXLqrl/WxDM7JLh4OZY9fkLayzV4SCBerIhKN7Lcu+pQxXjH3aiqx32d0UdIojx4
mFBvDPnzH9qDxHj2UJoREOezh90dJ63z5rsqz+JGCKf55XaWQ59tuP3cXK/mp7oPbKSv3w+xMFFS
EmzfYV+rJ+5gtM1ZvGNubmO7gZCC5U3c586Nzn1/2HsFCZk31Tw6dj3MHdlowLd6DoDNMOJ3/mPU
M7mo3nyQjLBsWXX+QxGFPmUZi1Xc1j4pXDG7tuKYZOeE0kzjlahzXlYSkNo7VljIulb507F83ty1
/WmNiEM9rzZ4d8TseUuQYITQFwu5AhVNumjs1Etacs5yGx3kw+xYmvzdOtM+w+Xls8LlpHaFQ+NM
u9KNfUpb+6QecmFFKhSF+dFigw6noRo+u9xqeKNnSYDH/NiU7tzxeShwiH3kdG42Gs+U+lJaEaPH
oVdJColYE6f5iSVMJfazoB1c7WdCGezEWHcj8tYMFkqnEnbuQy6lFYPzn+agHgcx3XCm+l2SSrtW
37bgjqhotRLrcv0k1NDTIoqkWai8PRbk7WUauzrdfHCaiYzA90av/xqehPP+p+82UGqFraxueHkR
xn41zfSTUvgt5r4jPO9sOwZaQP8r3+9FKGjCxYFWowTJNBpS1A/l4jO3SIAVBbhedd1/wZXzw/OP
3TW33Fc1K9AgCWOGfvKlG2YuRPAoeEXcoBwCommHdTtWGjo0dXlClAv91E7INq/Lcr5z0Vq/WGNf
E3tWCNI79IOBj7S0GWss5L/kuXoTI3wFgFRu/g2+bfsFvvqlW96MKFWJgV0jpdj5w7zvwDn21Jcd
h6ldTu4QnCz8mHXJ+2Q8JL5HZHtOEsB3c8i6EBhnkI6vVVfGTHyQvYA/kdxsMUsuxBqrMsImDfBc
Ly8ZvVpbRu4rCtIQoTzULx/KVEhPtsNZDd5loESNDGdTf1u++ma7DEuHk+J0UzJRiVsimsyTv1kY
/2UEB8mzd5lyoxBb7ubYTI+UaiMqBmnkUreAdNWAZONjlHG54+rljFLotePkb/6RNIohE8T4jg5e
qkKHz4B/XFxD+q3JcdWiwWgEwUcHDntBRRynFU2ZOE3aVHV6qJN8zrazrdeXx0TpcWKai34r7E/I
zASgO4DqqJGXzMjQDHx/9w2YnvnTvhx9UdY+zvlrisZgvM26nKb53kAT0zUl5i4KVjdDMhMch/Fj
wtUA+ta1WSwWCNm5gbnK7PpLBuHHh1muFVb2l6cQAcKMzOW+pdrKj7eSYFw+loVynJMS7Pi3Gvax
ivdexxTb0iypclKFAZikn94tETdrayDP/cY+0afATDMzmldcM6c3RFihJvUUNRhxwnplLJJdNPrN
6h77VZVq7Ce4keHc0/cqJ8BdsBJAc5CQb7bAun4UGl+MNDzjn3mz+EVNVU8YFjGj1MhVGBLZXBkG
n+epQkLE/czngmlgFzmHwAIY8a/NRTdxGkkOwuB1k2Vcj2SMFoN5CxQeeMB5mXJfAKwwfMtHzoId
51Y3BmtmEpbDUs2J7PcmY7kbrJdmrxAgAnFqNN7aRIn15HDrOJPqQkO/z6AQFQWcb31FXMIKFXTi
IRTjNVtyNHuKDZ7PwBCFmzMBC6z3agXocm1p01Q6DKqGmih+wpSRhnlY5hOnhjWJoG1eYr/R3Nyn
RKcOglmI3C1thqL5TraibiC+BBPFAYwhIApV2folIXcgn5/FZWkERvKZckfQKBr5RfrDuxKJm91U
v3lbgBjRwuI8/92H/4mSQaSS5Hc5WH7mqCs6qcZt7OHvSr0BmJjFn5aMA1jMVz0P8ZcsPCsbIhnM
gcON9DWK7D4rQWeu2mdXPAQKnkN4Qp8fdj2VLGupgy54NUNWGCM7J2TgF+HgnL3wy0VXd0vEgvmD
h0awz1Bak3IW3ptIzwRtuibUyggwk2kQFT4H/5EyLalD2T7sUMIS4hivgdytMhoPy7twmglpmYrR
xXdYmhlGTNmVCO4wIZIEi74EilgBwkZ/qAyYElP4+F5Fjl1Y8AXYZfAs9eRrGtbnStJF1PEEnu32
/2GMUER/fKCTX9fLZ5aROtBmrkAEm8q+FoIhb/zVdIfu3NP43gHg0Igc9kFzz/jwbSyQ9QtPSeYQ
eW/Fo7NrgP3xlTByQJVKKenqy5U/ul8BqMRqTHL6e9A+uBln912Dik0qbwtxpw3pj9cZkfuH3xCz
2VeNPDDkn87VRDF0/51Gs22u6QOLnJDf/4Ml2+UAfEN2ga6Fevea+Xbip+mT5WT34iXsvkkcpxwu
YvTCPqCR6pHSoFQjY6uloZu9RvI6Mnr7knHDwm7hIwqWv58ID2G6HkIecECoRKHQgaS6NPCDTfWM
LdIdIBfL1+ZU8zQuLgnyqMRnWyhVUBH+Jf+gUeEcBlE1ZShUbA0riGK5eMDq3Cq5hGJnzmncnJlz
y3kyiXDESx0anR7LNV3QVG9YBj1XvR/GjDE5FpYr1D3jJibGvJEJWv01hITs4y2+UcFSRL5yQ+IX
p9QeElJN5OE9J9gcRxqPj4uKhN1rmrSAY8g5dYILJNLQqlzV+5EUWCR6pfvdtTf/DxNd9euOJaM5
yqWoN9mco7Qz/s8gGh+esmhIXvLhSH0RkMSKhIhP/c2hjAvxjVevLA73jydE2XcuvnCAk6TcAfgi
KgN/bTSCj7aqBp9eDiDqLl+ah+Fz+MBHXG6JmqD8UgguvdMDQxGSBRHE9hqM0n7ceFjNzGNZMFBF
vIcCJNgY/w3+We5UchFTvCNYmDJaV8/bORRDnDy0LkphoAK3Hv/zZSVIEi/EQxISyqlezg1vV+vw
4WGNwbqXx8wIH7P7Kjoj+OZB3AV+VRfgXtrkONp2xKqAI/4CCfOZWeRXL4KIZlGeE6HFmfq+U17g
T2ymBMW/MfsDf9+Tq90nBs5o8UET3lgjXN+N+70fq1K52W7JsJTbNvbtaAhTRNB4/GKu5y07kJrB
XOrwnxH9PZSFeChdz+z9xos1whotSZlulaJiZHhhPJh4jg1d6teuosGcYTkUTNCycxEew6ayiNKe
lBB/90LRnsOO0SXi4zI4rpakca2kSncpxXqdjuGwaIKo3qh2rIs3mPUvgck2MpieM93dF9H2De8O
6TEWRaaJVOAt4UIFHAW8aaA2ocxJbL5H3bySwlSL4FN6MZQtr9obmIX3paac9XsV846m0KdTdjiK
8RRONMDKsP7S42/Zfh5ZCZvrMmXW2qfQVKj19PWZvTWnISuaDxIF7jNfYxGv1vJn9M9GRErb0ywc
zBI4+YNqTP+pWpkeDXjbCSv7YN4ALk4BFtJ+maHd1sHZGJLVFQFKY5pc+ADmWTwN2CqYPQvqc7WV
D3jGuxLFgerMIo0mVgThxUjXkHeWn0wwhQm7qVXmamT/itv7UCWTGW3tHx1NyhArk71aUOUWwBtu
VlywECpjTcgkEqcWRqQsaufFJ9Q5T8SavD3wJ7P3MyeCp0QlgTGNMHHaePlhXpbYt7wrhdOl9UDx
LAeYWiiMlroBM9wpJ4fbhkGYoCQm7Rg5r7wP6X8x0f1FCHAVsol4hO2ciF2v3XTJK9F0pohGnJ4Y
78jI7AtV+FHRv2J0878fcB1eq2tEN6KORo8qREbvYgKSJ1Go7AEbcRUrGeQzGxPSCrW/OZrQs+hf
FTi5F91KtAI28kaICe5RGkyusKU7YSOT1RerO7ds+ODaTxp8l30x9O1oTcA19oYSx3PhPb3BlSh3
QZsCrrinWQ/407pLZpZJ9k4pQBGxnBRsmIcde0sQJHYlxILwVKOyK7yMbxC6hGC004ewJ80vQLi5
d/GQAmRwQsy+4Q3QEhjDe+mXK9Pkf95c8OdF/guTTB3IeMItta4y020kTQwnhYaiiVT+yYsGL/0n
6YAAzb2q8QbaBWXH/u0WsjJM1OK4fynz/Uj0PwS+/djboRsSoeVqk4zc0MphChGQdBAtoGDgmwKc
hbDwBcas7mQMRkIX1M1JVYhufooHKOxd10vqaNtYAZpxPeY86zDGLixaf/7sX2OiQIttlemPoNjq
Gy0W+Xdfwp2xX3jlqTYEYUn69QA4YOBNlh2dBGB5ji0OamG9CZ8qLOBFBTkavswX/2OVgIi2unl2
CuAu4nqn3wKmT5HhjZeSw3NhTdXvJDrOEKPeKGjBmPQxpWl/RKqNBXGsZpM9ietNSw3xPMzqNu2g
zj9eiymOF4SNEcjVyv989DK4QKQX3K7xFM7fWDpcoC7RwiC9UIDgagb4kRm8v0liR8dXsRQ8Qqm7
egIX5rdTHgdnzL00Too3PFy1RY1yHZzwixo0lS74G18QvH5L9DxwD4feCYLNABpuWDKqFCPZCti+
awHU15fxwXpJP3wqOpJdFDBU+O51mtVdVeEU/+YWtIAZxTg8zl5uwprbnJs2vjm4aBx7QcJHVbtg
A4D1DdeNo/+PqcBdyKmNcLkCR7XMHe8I/zTu0tcAfZmtVxVniZ3YNY5tCNOotCpc7LfipOMMGLkz
wDcA2WkB+HgQ+CLdSc883D3M1dm3RgSnkf5iEpwks67UrDeXn9Ycy20WXN6KXKGFTCI2oqEZj6BP
GQ9ENx389xVAX5uL4HzDCF/fZwQkXPXG56S2jAy8PPB8iVG5KBfBr4TI5wHDp6CiCa8gCCuRoENA
zHyKNjqcuF1FcgkxnkZ3m2012AhOyS9LSO5MQsWHtDVb2xmA/nJnGD5E4xg7Mq4h1bHFyi8ggVWA
HuNaOHJadxWvaOKZcGZmj9gAPdDvyl3XXrgbUw+qNTnjneKSGeClblELCLmhmDuR3PxmzhogPr37
NrQ4DhXugzgUC+Q5+gFCgknZFM4JZ1/XLnIeXoh/5DIDjhp6DQi5M9FH4S2ocigZR5NLRsJ9fV5S
uF98NTBqozUM9xluBsoXB1g1d80VwalFKF9lLq5CDZ9MMd6xL94BRRX5HbPnn0zzDOvoBwnxB27T
79kYC46biCuNQGXMwK9zeIbD5Q+HpxyFwSkw68HXghSoMDUtOh3YL1jK/wLJmp31g4Pry0G2Guuu
y5Pfx198AoKGfFZKGnFGxC+ojeN6k2wX2/Jcy5dY8T0FZyngv/33sntdq5GhImfGAwJOUbbvxvSe
j0pBpPCHPcAE2qLL7RKLqUAgMrrp9nID1SUM+1FrI69ASgGGXzw/d+EYOa3jxf+1nSPHFlq6yhK/
OTD5gF34XV8rhAshQAxQucZhpPc9vv0++E+I4jCyuI0EX3p4+CyP10ySLTUsOx3mGaUvyyaed+US
85e5EV/Yr04t24Kl5f7vvvx6DV4sCIPY57cntio6K+bIJWo4bgvEBBSZW8EAONfwzDkOF36ki2OB
CKvZo9tmiDl18s5kpZEBrLffMsTUwLyvqgw3NSm824AQ08N2W4IWrcYBOmS4at1vbDGTtH7eN8ja
TXyoP0niy4nNHxN5+RwKbWL2vUV3EAC+zIunEhJEUWUgSP5dncUPfsHnddGAGXhgfmbDJzQ7Vh3M
28P2UFHwYO0V2TkVVyVwhvhAmc2vWMyqVrEOpAPgmd5He7Qj/fbRf+mF8r4OzWuym7GTGFXmTgn7
p6tCAjqyVThFBqgVoETCMVT1F+F5/FaXIdtRk3uUf+qu0SaqfJMGL8ZyYu/+8762tOLswePG1poa
ETux2LcI9G9KUbJkIJ9SN7kG0XBHo9+RsCbBYVuBr0artc6oryy/swaYWg3I1sVLCliPbCQzQKg5
5ZHxDL5VRgCxaRUUPuqULHhMwxgUBJFhdY6z5HCKmAB7IdFh/fq9aqvCOY7MTjtl/cEqleUWvEwK
94lqEN7BAzRrKj5NdwXATTGzZRjMB7EYd4fwb1KzVfDYWssI1QWwF2CHKOfdpkWUHlVWnr8m42Td
osCN9KB8uWQZQrnw7F5qXSGBBQR0G6yvHo9wSY9TOFbB8yV1GvsMttjKO2t/zE55MEcTADdB5X8c
boj6NUZUwRo7y0u7+Jb8DjGBuC3x/0dqKMo3J7ZmSPMo4K/2Aj4DFITIOL1jQd9mPmOGSm4t4lb8
b4iq0tqo0JvzzFDu/XeUhy3GPk0ijrRhk8okv+CBgdaHUg+QAwQ7KgUNo8m9yXAukPP8HD9Q8f92
snOvdf63ctWySwQVYQOLu22s6R5fY+WkDuWxFoeD8TAviFNoEeaC73L1p9UunoDEtaglwQSQQ+OM
IpKz3+AKlrz9IBWYw3YTEi6yj8rokPT6PCRuh9l0bts7XBFu2SHQLtZFP5e6PGWlc1+otPX2mDC3
O7kDitKiZ5pLCCTt7m+T3pGIw0wkTDkAdpnLvpitmx60N6X1KBnwDngBK/VGh9R9S435EK7+7swq
D8452z6aIwSrt0wI/1lkZX7eHaaeieAyoodNJsG/81wbCojmXJpz4YMNbEwPPH5NEnxMtpm8Q9Md
R3PLeSa5KBFWFaFsArJyK1P8q9a/UOAogC1qXpIY/yQ06yKNV+5wJqhuCvHgzPNbSuLM0BFID8uh
k/WZIRwVh7TCFVlSCahluaeQMKBYiX1xWOtAkhbCcDqWo7heg0glQ33QUiDKf0rVqFxV4YLly6W3
NVOEcIv24m4tnQfHh2kcl3OjeQL8yuDqNge4AA1RwIr/+qdnK4T/0FEXU84vOxKFp3wIcJyR9YrY
aN5+tPMGgMvYA8Ku/MENywGHQsVNzZUV1QfBQZ2f1Pd/eDO3JG8fuWUwJ9ztSV5augAoMUwUTRhY
AkD/5Des3gGUcLzNz32eA9+PtQ2d14N01HhKtPLdv6qH+/WNOBtgPF2UmJqtBqCkCB62T/SQVMop
loHedc6kNqRrrMEsIqoEsdB8SGa3v3Uv1m4mDgqbHZ/XBYEEN+H6nnoGGl2vagkyBC/GYLRLGhIs
E7tdphjHlBXFKoWFS5+iUexLoDJrlz/dyRF5uCnev+DAnJrBF97VQvRURJOhONlVCILzpbQFGyP/
FjywcFGkMYwtmIgdD8VFVvsZg1Ns1RaKgo61e3cChYAvjfRyfI3YE+2qCX3scXXk1I8/9/QsUJjm
xEKXfv9ZyS2/E3ves0U3hRC24qTaYiHJWhp/Jd5oAsrZfDcPiww9yiH+nTiwUuDeGUNts36iXmfR
x+nTRdAKbg/YSlGSKoXSIixku/76dVS3pZAi6mbz6Snv5leAjuK9VrwSds+/lOOcxlsBB1X2Q5oy
riQPaebz6QY7ERzkp08VIaL0wd+bXY6Fdk/K6ks/w2XEw+g1z/ukxVS8XdC0CVC6IxCKgf/IaAW+
fH3EPnqoVEvt5bxtT7S7OiBQ7exMdhTXmlZtF323EhBicUtfkf8xqqaLildZiCYF1VYo824RNR/5
8zpIuTOEgyoIIXyTBnxKjggSMgx3kgq/mwZoOrAg43Wp0o1t5LZka4mXi+A/RG12QHIOdM2nVbeK
zjuKOyvOv9vVhxlfku5uQKxxte8RwJkbJjMxZDsYC3/MCC4WlC9uJi/CV+jd7d+Rj16u+q0z3ATS
Y8Kd18lWgyFt7fi14Mx1O9j56bbNgUyO7A76xVyR7eICSQ5os/xB8iYdOYAbVpJqdY3qqWA5Tyqo
txj4Tfec2n32po+SSN7UlUxCx6t0aza3BGHwYYtuVl1UTvx5jT2PEUFhPhw5iw+qgAk/UCCtEUMG
3T2lbr2/wcAhx+5Fw2erGx3E4vfRGyDZpNAU9g1rMRL5zX9n7mYNSIjfa1pQpondnONgY+CuvQgv
+oNvdIS2FM0zNOzKMhs3/D7UICotJWTe2Hx3lMmDeENFWPy5qndBusd2+QlO+UKfhcWzMf21hmVQ
Qft7tI55SoHou2s6Dq8Gk2glS9glrLflENn712quKKUgadLpn0lMC9bm9vN+DY29tNr/zme+WRX1
acxkLheYIG0Nkh8zScFOD2OmxV1uScpMrknwMY0/GuFy01rIQhnpFGDaeMKhN5HdDgpIGiE/joAw
5YvUCC/pR65xI5dFys+pvVd8itBdo9eM1sm/g73X8lsv+0bgrEZ6VGHo0BGxvUOYyJGSB8f7hc+d
aAHtF/YPkktLi6qlUa0bZDtr4nIgDALrHPmwAQLwc4sRNmbuaIrvh1qyx9JfP82K0iWQIvxniOBn
HN06n+PODcXpNOL6jB9rVeglG2de3yjXj20JzAEp4CkyYL0T4u60KbE9N0rL4JHkEmuzMo/rcgAK
wi2yPOs6bgJNTZP8Lzj0ULqE97JrwfoaZ1jt8mvTHmx+rl0pXEUhSFsm/jtWWCp//zsaGJzXy83l
ELehliWfNjBWeaKflsuGEQVEZlyyKC/7Gvbk8/XXSzcl/+t5s29nPuW601JMzyaNTb9HiXpvgH0t
WA7P/BWN63wp7wboqDXHo2g85UraDJ2NPmhx1qglgLiM/vMOvRFrKSlDz5eV7DDyPcCpJnL+Nio7
jjPpdySOI4GaVnUBMRkdKH0gNcOIAp+U2WI13QwgdWUkw7z/JS57aSLMpSwz0YYpd4bJtSXJEKFw
aMeoxE59GBEi2b2xIqmKJch64xrRmRrNIGOBwUJSEoosip8dX2oK3k1hO/8Og7qHB3GxPaT+paAj
xCql21XJoB0lCbtB+4z3TkS9PyLsj8fe39k5fOHmWS42GhJda7iZ4XufHbEAXJyLCAaNz1ResuS3
/i1nMJVrk6IiWEdsTv8iNyBy74oZmp1czdGuP3HJtlikQRhgLSeNAPathNgi1fabjNXLcRAQhMkC
s3p2U4fvqfAJy/qigW0QJQ0TuIyYdwkerBi3grltwqj/6H3vxg7g/JHOzFoPluOH0AFqpDFCY8SZ
h0yV9cg/Cx/TMZYMT0hy9B6zp0FtwipvC8ZuzO+U7iKGHeVqYywo4RgAkQ+oahIL+mpRkWtn+tc/
JpF+nCWc/hk0nGYQvQtmV6XpGPGViJUtC5j6MxaBqheZmZzu3PQ+0e+bH89Af3dG94Ri7BO6M8J1
T0RHKfzcUMeA11j/byTO/NSH2GFlcPmySTlLogRLJ6K+D4czMMKsSiVYPb4V+6klCIIlQzCjz03k
Y5+5LEwAARv5MZu+srfziedf9OV8xRDX7CES53w+nixWVDqCcDFS9O9xCH0egTZ4N2Ycqi43WGhd
AGCFqWayAI4i+6vRzv75zjLtlv2uuk96cykZYn8XxRkGSN9QQAO2jM7mwT16GRHS3cLfJgXRS7aM
VPxoEE8qwuxg/tMo0Xud6aCk2VsLk6NphiqKC5ZJq3/SZwcSgFuizVQeY7EN0CNaN+zHIGk4uEWT
e7CJ8TIledrbP8lesyi5g6KeKdUuW7PgGQQ8stIegWmIFtwjuFDuSi71/f0b/9tZVAbG6KFpDAzF
a2v4H0DrFw2e9JGYe1NbJvxQqiDQVBb4i0aEWZnM7RHKcCJOoZvAYeZMsCpeqsAm4Ke31t5QiJon
X2PoWFJAmW9k+qRKYRHMqVMbaoFrluYYTaRdeTxCU15y1+f0/BVWrU/F50C0AtC7rnapNTOlDBC+
BK6mbiTM/Uxv3hlNZywyyVCloH8Kn3uVE1wgnyi+RawtLz0KP7US2vmKfWY378UCtvT4PcvDycMa
7XlB0haG1kP0gj1L85KQDlxuI5PGiOQswxcQ35ju3fcvQu+ampx4LCmAMTLwgcBPbs3YI0nNLWZc
4jYnxGiaZqYNcginYlsLspe3nZobsEndI9MSJjrWkzhM1sfYSuYoMDRQFmuVxc/2HCrIDn2lYgbW
4F6BGHuYQb/94/AM5nCpe42SG9hW5gM56exQCtukeBeDoSYJLvTzFNw1cLpPQCkJWtybsYU0oHS4
Q1ma45YpjXnY5W5Otm87EfidJHetvokmKPaQy4edT/uFeMVjVcR3PlDNB5Wgd+NlR3BSlTeLk9Jj
JafSKnAxWTLZBsncE5xY2tbIuF7CjxkSij1F59wVah6wLaU3tVG+nvEdSlxBhiPoOVoCaZqSdnvN
JUJcuPN60YaUFroy5+SCkxtQHXv5tXMogGa4WLz8IjJ5AI1LxVZnfpVCBe8vxotxcQoSs2yNQsI8
oxCdOOChJMsy1ZO2nJQPz3MxUAQS1KAy10tO4/G/xsDLlVDNBFieCb2Y8LgWjA9DZN3c0BefEPD3
iO6rsB6I3PbF1sOF37VUosx1JashyV9EvxbAu8kG4OdYHnA8c0LTNsubkVnAN9GTP7PsCcP8srAr
8H9Me0mlvYi9exGx+vy44gThDj6ftKJ7n0i1I1msONLrdFQr3QtDmAq37D/vPaqUFJ0zJ4igdfL3
oLPVsEt6HtKNfFByIcGvdOIdPFxYOejYfKDCzfC/IVioFTlqs8tZ0F9zxXYrbfaNVEuMgtJPxanI
m3q5T9ObugofGGverKEWs3Z6VDQLySHH0rjSBMHcu7FDOnCz+WmDoFdn31TPNN2R5vDdJ0mN2ii9
tQDr7tl/QrOqoXRPZ+9O11OYp7jGwCHEQRupzcucUEwRBCdwyWm+GHMcxAGA4WuATP9BWJCrUfc6
CH8kflBPNxPsHdGQVKfBogGZ6uQ9XGaLEBMcV8+3v8RHhPjh0kqtLJVSwRrBMK+TC6HhIYj538Qn
hYXVK5oqmYvDKNKBRq5MUq7kSKcsipwLIPmqqqVVR6V0/yzoGLsjjQW4dtaEuei7A2172/ThPiy7
0FZN71fa04rkQOPs9uVX5Ptl8ReyCoUo74dL378F5eeQbhAb9wDzqZ3DraGWRwRNl1VzVfyNZXv4
ggdGTXz14FmViZBKqd8cYyfbRGUgdWoEqDyicnhpMkOKeaLA9x7WfPiGEOYLoOLeyUc1PTjvo85k
P3Fp/V/5Tjty5Rncw80OfqEDUGQCUfOld+bUvvKe3Nb5VSPghPBT8KIkOJQcKh07qkA6SdsscOBB
3HxNJWG9FIHApKtKhff3EFwFWcU5iTFIoccPNppCR0RO1c4csBHYvn1y0fvIqu5UJO/fIMDaKD5M
DL+wfSiC9SmYWHSv6rG/EUikgvQlm0RNSwqlNHaf/SL0BIP4XqfSF4c1meuEVThe84KL2OS+eJXM
p3uRSFk0OWyflFYGyhwIPmMpuvXW5KD56tjm6tExX0ySlawZcT/I5MSVnnDZ5wKv9nT4kpzMbpwJ
VPiRX4K9fk0KN6ysr+0J8JyhyHRsKFfgv/w+k8TKQTYP8u9NaeQT4vXc73Xmu6tpXmYFPApwmxar
nMrWseBgKCWk68C85JJ/QCA44Xpx+7655e0mYKGk9iF5MwsBY6k3akpbQ+9uhk74fSgrlV8O7mZf
iELwAFK6hWI4+Jjm2thnqg31vdTLRYeYiBJIUrM/foTMDr6qvEdA+hZ8gXKHRDF8sN3v3rshGw7h
VnfLSZD/C6UOIi6VRVNBcl9fJzuX5hjkvumuJuSgggJ8WS4iaN5FEC5VCQvv8XuZc97cZjqWGhWF
3zfKlJ0D2hlb0P5UGBu17A+ZonKiGxHwJ20QTuD5/6uOynDMDGZdIGidRYr0mbcnR2+sn06QoN28
RvdYP68qOcL+E+pwk2qGyd1or9+3t6z7wCyJkrOS+J03qKu6BbP+hlEdAW8Wnqf1xe4odIBfp7+W
cIb2ecRKdzqxNyIz+o1ybKEBLHk2iw1v5Ut2zzWeeOXBLqkmKZypkAWWK8FB4x+7uhMEeI8550Zf
gd4RfYJEsEQ7BYHtHNX7LSJYyLw5UDsavkJfw0dii2RyVS+ei1xlZ131VQvA4UPgJ0XcACTfGO1Q
Y7Nm1uDgRJRFyQ77zuNcI7nxqm5Hmbb0UhWV00h15bnsIcXqUS9KQVGeSDKdjDNXEyeeUmiFOG3/
lWkzf0+sRDi3XZEPzXhIvIwHmknLq4seIuQz7IrNM26leiACE0wZh8cGRXgRPCsZpyW81GwtLP72
UypEmjZmp0dP+AYke3anB0Rl02PgleUcCsqMXunRzeevSegI4/Qa62kVYu/F7lQCNhjEgd0fabIg
SL6pCMXi/XTK6yacCrejBM/vK9UdOCr2BALcSWQYbOwV4ot1ignmqiBnp3btd6VizNNpk+5JLMeI
GeQ4JHMr2Dtc9biX0d+qK4+HoRTVtmbVD03VkRTtKYTBeqQ6fXkIoT8qb4CPtn89mmvGU8q1+Wu9
LYyW6ts91Dz/Of45ZqwEryW2FhBLQSh7UijOa9guOkTFSV7RUmBH1CzlXAEDbrEydVcHuStj39PW
rowmFi3M2wc4J9UxZq9blTaXYXAldmxXPVeAGsiPfVCyvVitoBkJpJ1DpCbcEhm0j7m9lwQUJS2a
CscHxWQb2Fk3Iz5u60OTcEAME3ZAN4hzL12cS+kOM3JerrEflN2GSE3OffQcbsiG6foQZ1/kqLFz
Yi8tk9liFOeTAS5gxBuO5d6lkUSrWXHUcBdRvPdLCko5jcEqO37VpK3esHVxoe0EH4yCdynqwL1E
VYdrgE9YY8Ej7jF0qlNLSeLmBPZsY23vZTdtIHcKWf1ZgvRVKFr7xUILqHgSY7mGRU/q80RPZOdn
5Y1jHYEavtt3WywFpWp5f/Zc6hJ9g1AQ+HVb7H3PzmX5kfhPH9IAUXv6Agtx9JMFMv6D8yTejfWt
Ql83Tk594n/on26DEL/H1QSoP/qi1ft0d+YeRXrX1/R/kxnNcq/HTmMMNhFUSR0B7aywacY8lvUV
hmm5qhIMiTptT7hXRboggNbirf4ae2C1FRz8nZ1Aqlshwr1A+uvG5UA6Xz2icyvC9R1i4OnbuXdH
6x4/7obsfa3Ya9KgkilCQUzv3MoJAWUygDyOwvXw08hdsUyC3iZmTPZ5NSpRUsDTMg340NqoTGFz
ULwiQkKSGyZ/B8kKSS4y2sQ3TiQ4VU9Zn9v69v/D6KIRCnLB+TylRjOmLOicEbkp1q3r7czLKiBR
y68gPsrilSBY/W2e9WKAIQDQEntD8PYTTtoHeRHGJMDjhTNVyFxXGSNFfvNazS+JmQYaVTpsI5jg
Quv1J9V2FXqunWqYR8oc29nhvCLNiHZG8+URx+WARgkyk1RGd2ztezdVeW5mudqXSYxTCcfBqB6f
T1TDqSKc7SX4W+3nkbAF7m71Z4rQB9hnUg6FMUjr28K/fkvnnJlIy1G7CCPTduAXOJke1BZxOeCO
fSqa0SHuyCdLh5GnvSmf6FmCHU0LQ0Mze1OYBkBGW8mAyz4m+svvcOnZvskFQolzrWxrjJBEiFqJ
ZVpdKD6NYOWdSnitns0r8s4HnRMn7xBmtjKfa7UX67E8IOYjdwRlWOz1dOKZwn/BY1ipTZHsJYzv
pvSjBE5I+39UyUYt88XkqoTde8dHietNG+QWbO60yLNIphGyAcjGPgxXJnxi6GOwfiE5lT9P6mXR
QO+AYbjCWCpGSN5u9G6i+GtoFD1BoUGWBAq2JerW1aJ03G3+T0Cn45vVzHu9mWfIuKa0Y8ZoBGcN
WIpRzQf5JGoYctZVAcyQMem23z08IYWYcAfLiFh0BSK85sNyg0rd3gt57eiC4fBDa1Nw2enwLKA2
Ensw/huwG6J00fTKhJ/vgB70GM6MCUIWzbeP+zzh8lakvQ24Lyq3jLgQF8KbULfOaLFixCEBD3wu
0U1bdCOnuZq38qDHWIDHJX8Xh8hi90mXM7OrOxUgwvyiSYUg8UzEIdBNlURcB6xRW/5hK6jf8E8+
pyn+FKzlwHcmuz1y+UG4jKV2k15HlUfGGolr/lbRh4BhXhpVIRFxOf75sdwGUoNgnt3jUgQDiGhc
vYrDiwI8c+OA7PllVUuV4KyJO5s84U7fX72SoEhSuxDPRy/RNHjtssQYxTtU367IOSbScQcEn/85
ZKMukZiNz2TlBZG5APjUtyiaxZewpm6UqprVhutaGQR13uSXxvPh5lqfLavZT1/WcNeiNA0Y/9Gl
Qp36nwDm7gx80JJazh+Rz3gwkfMpBMjrxEToWMAo3OCUttlkXFWrV81KXzckbUZgOo7OKzsElQiL
kqUv63T//RkW4k39HHK4vitcOmI6d44L0+aW/GeKyViB6G87Ha3qrKNR8j2sQ2E8H+Xrhj1DW8Ap
lCfcaHKmR9jFoDmFR7V6IwKyC2gnhJ3sZ/634ZY08NYpcK3rxCSDRyJNbhfakgQBGNnx5Q+/munZ
v3FiJ3m3E3KqhowPVwb2+8W/wnAZHZR2Z+UwHCPV2oZCln2zD/Fc685er3VTGEiUiOCH3aygKL3i
eGMh9/GMj/MWBCcV5a0VYrEGu/1xKre3FHN+gwp9xhIjcFNDWVim5x7lMk2VarCX9zndYkXahgcC
GPpZTlEWxXyG7l84iPNaLkdcdKd0ty4oYjZuQJxSI7uAkiOKDgIWgfLzbvYWGaQOYeOd0xuuJy+u
i+KOxRhVOi8T0CoSZDXRQFmT0uke+q34+Pu6i+jGBC2h1de6/G0be5PhRVCqiAclguDl78CjhGoB
Z/N9LHANTdoJ0Ce9B0uDDUEZaIt7IjG1i9rkx+ORxriYhawi1u9IghPDjMxKptTmV7egp01Shebv
zaVsWIzJUEUcEJTcNcXB1p4zcJiTBZho/M1jaboWi+XhAHHTD7QWryFexzoPlCaXZPsmgC5DvWD1
jYhzR8wIL4vpXcMzIB7nKUB3NrAq3+pjj0keKjuPCQRUq7hRl5ePlS3ddgPCoXtf/HnRKsB0ktut
QQjJUHl/8PU3m8MQSccZYHkvV5hlItqKg37V9M7UxQkbStOdsEUm9OeLVPwBMiEpTFrnnW/PW8Kz
BoD6ff6UHAd3CNl4j6umGrg54486TCnRznPEqJLm+t4rvfBfPmp55KakIl3pZn2NRxo9DaIJx64z
aQbvBtw7UQw662mekPu+fd9aZ2M7KEB97+HuzBoGAkjdyrs6sxim/7oS+nnIOrnCPVpxkCZoSK+B
/4+0Gag8V0KxfbmVjkOmik29QuCzNuacGnAu8oTU6RA88Bg5yqIeKNUlZJXe6Vj93NavW7SeX6LK
GYoZ2BuHGWuD0Zbagc6nTwJJ/smIz0QNWQWB4H3UrmO23rNKqaj8UaAOTmZdJWl5fQx5kGbFfdRt
Kc28/VbtnooQfbi6AxNMIP7rhDJpz5P/XHGZtRQlnHLO3wDGMbOkMlZWtG4RIxBL/7Qkfs83xIBZ
0y/CsUOnQ15GDhUHFNTYJBA3ecA7CetQFYH9GUjKW3GJ9zTdGDFVEMqXvdV6nsoI8L9wz6q7tPT7
+4fQ1yYzkoqs94fHaCZAfBF1U5FFiI+1rFWxUTOa1edhDYXsSGAfiA2CfA9O2KLhQ8eVC4BdPYhJ
eBzN7tjHSKoVaLRxXgpT4BRBFesh16SjtkSqB6GP//1ymuMqggzXy4i0P4vEsC3D1G8rU6TH6vBC
ZKXtlkwpOhicjUi8ExPehtFWB9taZJ3yx6yDPq4iygsxDdRs0kdrksCCM8omgg9X1V7fQfll4CBJ
BbmNbLRBttZ8CiJrAqUKCnbMWa9l/A5rngDyatAk3X20OXYHdBpl+dsO2vKpuRWupbD734dGkq6O
oTf7uhuqxVUz8IVLkGgBU2+mWb9AVF5ZUWDoQP7DS5U2099voST1IkgcX01rczCGA6b/doV3NuWE
sD592dxaUbsifMUHcpoJmZ0jDaeW1vl2azRlW2jDcSuXitsMVcICmvG/NpHUriZ95Y9JjO+D4mDO
hYTkXdrQPkfhy3UYEYGG8I/121SZqZFNdKaxMWwYIaui822POnZfwf589DJcA+kXrJSXsq//KKkE
z9qvObil7O4BAN9UNPWqf1mxxddsU2e+w8MzhXwQlzpVnFYEUQ5CggHQgZdaqYE/kHFhvcCVKn8r
G9wgTjAnkg5FDniZCZvq8/ch0+5wGs3cqx6zS3aqBDaru12yNVDz0LiY1tyEdFqrTve5C2kzJdM0
gF8P1ATab+1T9KCmDVlY4IhOC5lgey5RLTl/WkrW0lEeixcJYQ0/GBgkntwWdQN43wpOlrHlr2YQ
rfeXODQSpjH3eTUqQZdr5frSR3AD6mxzIvt5SSQqaBrbQsDDbHqPrIlZdmq1cbaA86hOq9E9ggio
Wkpu7GgVnT3wVNU/44x7qCfDI7+FyZYjNJGAVNxtvqER3nO2rADGWvTcB9THmsrg+yNALV5e5gPL
8rvsb6uj/gLro6lFZjFkgyDcBtOzdffSy5O1KgFNiK501R+kQbFcOgr4sHrP+DEaeTbQFLbNgTfk
+Xve0Y66hhGS7+KasTlWLab3UiK7mpiE9aH429+k6emVTuj8sH51zfO54qxdaqprKnPlxI688fjJ
3E4zjwHLrKYylISF4zq5YAfhyvBoCMwhJ9gRys7RBYuNM18taby+n+4M0JOnEsOdKLDGJ1qk2vtU
wuSL5aCq4nKlvUupQENZbEqe8jFNlbBl7W0ODpaLmpEEAtHY/q/AeHmkeQLQ2uJRZPpk+l1p8smy
VpImD0jpezqtztx5uQEdew7SydhN7Isq/P01FQPYSIGr1m/GF64G/FpJwYQJk1t1708XOYNuQYga
VjHZKOVqzROxY/bApfnwV4EdEvmEfSyN+VM/elZMkBu1ZV7p9s2zoavkaOQD/xBQYK2BRwDdoL5y
CTBZZI/y0eSss+Ck6oRPPQUiipp68g0PPV539Wbc60Ia2gfb0a5DWtKF3J2o4HhEvvnOloCD3uWR
p/bNsmBIhlmuDzSKDAipv3sYvFaccw5yPES/t5ufPQ2LXaWSGKrq401iku5ISMQavD0igqF2kEeX
OdqLIOpVcgySr07DW3/nMZmrowRHANcXE5gumXu50LObJpffisZYE9HOi95V43RLt53U58EUwSrf
u+u/nMMm1oJG9zRNTJPY8/e/383sik4wEVrZYWa2xR8dxshMxF5mlC7oV63WwHpsIC3+e13mKNLm
UPzSAdj03eWMN3s5G009e9jkFf9s62pQgEoWxsq1b8tlJp731hEJ4mcz+qA7dso5t2tChqs7sXy1
0PcBP7KdrTHCM+Veox/dh9ZQUn8fn0NPYPoncHMeHHlwhHWOOXetLTcAuUm/UlBV3l0HZ9oE8EFa
uqS951gEwu2d/g7qOWACDs2KMgqvEAhbyIG5PU7GnkqqjdLMJlK6eXNAWYLRRa7DTyS5/OYvRYa0
C6/tjLFydlvSPo3zLabnpwq6fq5/qpsYIhfi2uk6o/WItMBN+p81kZJu13o4uP4Rzi2EZxSg+ubU
8WcmFFvbgK6x6uOXhMtFXvRiY0uqxwKNg1IF5MnL15hi9jqzZpe+KbxFomTrGx/0LlAJeuDzgyBv
Ixj1+1/M1SpCuWnnZxk7QG5punCQVSKewW+PpRoxmzpfrmaLHL9U7oPjkZ3AoXZ7lu8JLqR8UxGj
trgVLXRis7iydMreVuWFKCstDNh5D7B306KxlvTLQc80VHwl3PfmkFaGs59Q0z2reKqaAarMgEj/
5YGYLnJyy5D8k4N7wyBDRskGROvdv6JavgZL5bsZo1kfCushkLXUpzGGaJrZRhodWqJpDFRYi4Go
0rPA7O1IpwhZKMlF3BcHU3EMoR2ilvt5Lin2u87La0UqhUTgz1Rx1sfbFZWP4/nR6kiQAy7xUxDy
oYRtHmniKyVy0vO2MfsZaQKye0fBJ41sN1gbHc8FsXGU4Fo8peS2eF8lcxvI+h6aPr5GXFeyi9PH
eGTlX62dpjaeYr1/Xca35O6hxGmGxudMc/GH6nmxzX/WbGwxfs7Ro2DpEQolVEgpn8apBGV2KS3Z
h3u2A6mevABcbdJg+6lZ1Yl6r9xF7nYf0JiVYcgZ+3Vnb9SGwGA19O3wh0A9kzwXKcKHRQQiy76d
T1d/DrI3+EBV8tMwxNdlRpHYXwAPTd6irFf0La+QzVUITpLtKydal6puLe0mZXwxsiJOKmsL7tJ6
DmLyYWrRD936VxXLIsQr6nSzp+pG3Mk4nzJDdm+Q7H63SPxVgPi8nn9NMwpBRfMQULSYPjLt6ni+
8Gcex/KJSlTjKCK80Jl804WLnrrxJb7lt5Xwudp8Rij3N2LJV0yu0/O/2yEuxd5TmuEbl6oBsf7K
FGANISYRNpXSm9w2X5krvWbYlZudXdZ2Azchn978hvsKv6ZVYBqzDxowgRt+xSVVPlsDjcrXntH+
zMaAOTFh8ZJBLZ6wjzfms7PBUZe9InFG1Q/68itKxq9Et5C0SEfTU401hWlu2aut8/vxc/XYLAi/
mbJH9FJzSp38nynGsqSslFeT/BXOJPFa8Qbat7pDNyqGE6Ygi98L7IIZbV4lIA3UoTCtkrVM0yOM
K8kKCGFqnoTkCALWeIN96KSbOuY6EIrVUyozbLuSOrCwPyykRk4IdGWjh1vnOnG3IUe/1SNm5inj
N6SykLguokOWeukXEnNYgzG+gnpeSqE5nA21Xig2OeudE9KLZGCQxycBtNsU9ZLRbqK38Pb0AM00
0lT80llwwE9RoX9JLpK95Io7DeQRbejxdTgvCRU3GmahKC2nRokMHih3N0B5rhnJur0oPwrgp1UB
W6eIYDPnr+/wgUxIFse2xK4LAsxbNq7HKjakcn4c6O4TNAC+tjDJDqvbXzcqa5dlY8xfjX7wOl1y
ins/B7TdSStoEtnJolSD5xn/SS68cpBE+S9k2VosStSKgqzVNmENzGcIdDgj7T+KwsT3ClhRlbAm
Jxun+Ry0IDe/gfxN0VnqrrLBpcuORTPvEVXC1nql7opPaHce6H+Yx4x3f5bnSJbakLZi8YS2CO3r
Hy9NBflWrTKY0WRuyCjmd8EM2lmJPoAeBdKH8lx8SXQ49mbcGYJW3io55990wK8OzKJiLz1w/2Ur
57dbo5Wm8aHdhHXrDuKb7grdcJ2E3ZN/FipJMXbNTPkbrLbXdSGl1mSB7EdJmFa0thrs6wCQX73d
POWyJh06dDJ1Q68ptLadLYNC+LQckNaC8Ms4OIxpW/ZzSuubKQZP1VDbOn0DKritAl7zEk0meZ5E
66i3LVla+g6HwEwCCtg9YLzTdwCM4m166XcsxY9ttXYXt4w4aXcoorrpWCOv3C3b3xoww26Oa0cm
fhRtQw+ndlXZWGU+eCVo55X2jKKWyJ54nDcBLlt0GUOV0wEkts0oULip2xnziz3eK2Oyx8WU6KaC
WqVoUQJRxt4KZr2WzNkLJ57LaHM7FVUBMFocbxeI9JUA0HnxY7n9t/9mzJ0ZcVFMQ71TWmvs7VYO
JGQ58xumqRMFABJhGpmKw1JUXGNKVyZB3j4oj2mHfnIRuXO5mFNsNt1LECLDYEMU1OXCY2UYcNrm
iDqa2XBzOyD9IWkitUaPhbx2bzzvv/V5yx/Yehjd3295Q+P4843qcyedqP4sJIfXzQzT4etdYO+J
OWH3ghE/Qy5x8sGr4MktliyvRGndWnQHG1Swz4lze2MBWbaBSD02hhYqMp8lSihHxJTELtoEeSX6
Uau/c0VvcdGM9MIpAMLgyEkcWSPSyGMhzy/HL62SHXwcCPZNv3QwcWbcTjlXLzcivwXBYIocoDSO
q9AMrriDn+Z9cnJlPoOvLUpTYxLIjcV9HS1za0Z7J0ZFAFPTh8gPAZKHYdgxOlTzeqwgdCEBoALG
PfMCcWhAsSF8FrK0SIRpwx2ND8kmNUpEdsNolxki+X+RSGzmtxIkRU8mESiggHw7xO8gSGKDiJOu
Pw0o3WdarFT6f1rVAD1NAkFrfJtJ5n9Niq9cEbiyE1wNZmgo0tyK4Ot0VaUsBv0iVbjr4d/zpz/s
riESHi9jDUIWiInwjHoF0TinBDGEO4QFLEd9WiNUnbqMebSFc14IehvoRO4h60QmrmzjkolLMhE4
ntlyyBK47FONDeTMVddMcGfs78BNChenqom2c3Hxxx2nFmNh8TVWU4IMupyvwr8/hUEXVc752MqK
tzVArR7tDUnA6MfrQz3XvXA0hQYzSUypolQh42Nu3+XwVw+pzrlnJGlrplcxAZtzcKDeA/nUsS6o
7O/mPfxe1vtDZzKvVl2CK2Uym8JJLax8T9AzsWh6qGhkvR7PFux94M3V+SoEf2Ws96cNMBcKzAb9
YfuUWNLqWd8XdyswHUfE5h4k6ovnVyKVdzY1oN4VeTyTK//j4Vl5G/Jc1v30VTw8f8goLT4Atx/a
fUJw8jCJx7OOgXrCgL1Vejznx4T61irnyUuZ3EwBUEi5ksh5ROKN1QvewhmFCQ2ZczHrpeHOTGZp
GfJb5Y5fzEo5abm3toBwDNX3W/zvh5rGGZ7Lwtkhx1puzUGooUZhHYg6v22GFS49VShC3Ofpk/f2
BOe6fJQ9DwJUprBkei+xce15x0sR7TwvQf4F+U9WyjY1erDXu6p90SehCqadL2s8F4zOpXiET2RD
0r0ZVjFUmIoh4GfJOgLDsmE7lZR4lqiFkyMG6i390q4K89TtZ8hWiZOaf4iqB5NjNfwiZSzRxC0X
/oOtblKgaToQr2tywd/9PYzrhOfD2/FCWBU3btKzrxjwurTmeLUE5aNyBrg44u6+pb9agi3nETmZ
J2nXXKwH4ceS/2FrVm2Us7el99/k4uGBvEz9EMyNyNT370mX7U4Q3afGXM4+yHfLIAidb9RdBEqK
S30bqb5zQsbbIsskADYav8FJ3xq5PCE8A4RW43d3kwpuhPhtVG2oXdT3aYAQWJAQwgRocWb7z6ed
03ZCwb2Gq7ZPfYXvAlphCz2YDSTTF1fPbsIP09U6BsEMgs3dcQp/VjgahuseKvAwze7TOGBXRjvv
X1M83lFILyROCWVg+FSKrWc5IuCCkT5bKjTAt02wNE0sL318Cx+UxVxVHfXfdT4+BRCF+4YGmmj2
dxR2jp0e/9f0Ru2mGIMcgsVPZSDOVkAIg4enz2HWHIwCmTK56fRZ/xaywefUfXD+PTImk1QDnVgB
OL4OiOBifALackqUJEWpEBoJ2PKAMpNKUszOp7niKZp4PwkBlsv73iYVOoyfHg2yJfV90vEndlom
YKZl/8PRczotGZnNrZ5np1ttUAEOZZlNvUxNLpWawF1g+cdgyLvOBqSohihs0VPf7IT+aoM220oB
dQtnC0szYpuXfAzRDb0D+wkSmolOZT53ztqrY2ZAXyQS7vRFF3Chmo67kynI8XL33qgpNWAvby+W
78oRNicPNt9BmvQdPaLrd5dBW+H3MGGvGQ22jvqkzTuGKrkNgA66T0LHxem9Gcb8+h/A75uUGILy
XKcSzIAgiFsX84Bv3bAYpCii6L0nTb4Aww/FfkHbw70fv6JM1i0MPwqCvGeaspe5e5rB63Pbi//z
cFvt7+2VuoyhMbtEDs0sTw+Z7L/qH/LgOtpXNxHxASxbOHhPj+96zszBHLmLuXGm7gfOrZjxhTRI
H8XuY7+503z58bwZK8KbSziWYsI15Kf0CC5labIGc8zCAU16z+cSZzkBfL7ZWbZfcOdjHS/4Kd4p
2AI96izKPqnuHLI+FN6mUZ5E6nuFzIZbktQOsw73Lsxro8RyzsnHQiT/H2wzigm1UC59Di8rsX1A
OJvgWVJaAIEH3N+mRuLfHFst60N89VU1hqty/nSvtO7SgFDODlFdAtbGtYdbBsUBtOsEXB78BGhr
xG8EhInUua/dYZnqWZXNdfrLsqr4Ok62/ipfWeqt+mdxBF8ElDE6CbABvggxALG2DU90DM64ePh3
rkO/CsvryAJsdJ6sjnJ0UvAyQ3l6t7izynFCThDtvnQB70A9HXsmIeX5Szkqoebx2FjD5LgbYVwY
goX9Psq3siC1TgdAoKsNsdOBHAJ3dOqGuMC9ZfG+l1GqUCh1NRJSOiWmNhW/whDidBhKYdNxJWUV
++9R9Z1Gm49mvWqUdPu4K1k9oSYrYYz9+OaloqCBimVyKIYL/ppu8Dsl5TgjGPehBJ+VSO0aPLiy
b3yqGxwtuwVbaMUhCNXQocqo0VBn6xhhrfcmVcl1HGY1dfrmJppgHakQCsO0g7NBHxQdZQ+FESOe
HhdFaHKJ8zynx6EtziuV7GTn/3KFY68/b5uxk0kJ9iP1kjGC40nBsrzEf0lgBNljT4cX0eO6f4Ib
yx0RSawob0Jh3ffYfSf1gcUvnHsNm/36WfU61yb7W1gBv3x8ZhkE4MsYhuH/1bST1k1IS+z0ZL4r
XDvVq/myyrdyvWWrS2/+yX+4dinspEmleFbhvRlsnoXn/Z4nfgTivrTaGvGWD1ABlZnSI8cqvAWv
HqEA0S13WzKPgKvge83iAsoSukcG6eMFOIGbxUE/Spaqhh9SP4ZLA3yj5sEbigDI2lTpVcKGZKrv
5heohwlZtkm1AnKfhddlGvKr6FuxZ2vu6LojpivdWNVGZ3kG3aqkndnKXPUiosQhV8aLiL549ib2
ZjD+4B2jR6biVPh0wIwyTrV6JsJB5tsEqKNEOVl8NtPPI31AdaZ+6XCpbtv+TDxuQJwqgBCEUXHk
7PvwT6lF2pe3SnlkjodtQ3vaGKVfAIizt2hIBV/WkEDlTtF9CKUO8BsfXuRTRADWkyzjiimc0pkN
vjl0nTQTlQxhnCEPIHXNVavfjxlod0XhncX1n8AgkEyTAsDaI5HutDB26jrQMXhqCiSmhnTp7dHP
P1OeGurcPMVgMMBX6HnYimIF+s8FHHzspYlRJ7EIvmkOvFb2mlTd/M7afJf+BVAaTea6WLyhIqSW
qeokbEazlYRyI9km+T2d8iulCjaW7jV+BWQdboNmqDa0/BVeHN8eAsYPJlzrAjr+ot+MLMV6zIml
7TdeOzh1d9roiiq34K41e+PzJvUFpDxCkomJagkOk9CyAhh2r2MWw7PNPEcLqx4zPGnvUye8/K/l
Xo3xy/J11XYI0wiQCDA3p+EKDWamJNIQky7gtn/srOBTaxf6lzZt22medqR+mjM26RiMt+4gsffK
v4VPX6VqGGY0pWTEEHNNI3K+PFbFdE28qTvyGMaS9VLsEv0rZj7b254LBSrtfzgYciJ/ibQfGQeq
2yowitanPXh6WA1lA6waFcAFt7u+lBg6sMbUZqo9NgtitKLCwRNdB05Hg8kEMHVjHA79IJb7nDBh
mO/ASjhhBeMPaCwQcBB4k00xYjnw12ZPMghr8DdoFKt/wKVBzL2qu8v9qhIV4Tj1oaVYaQuJTaQ+
7fEkZtD9lUYk1cN08Fe2n+cuKJeYKpixmcMk1NTY9Xkxe2Fzh0kylqNBvECcPU3cIrZ13LorO2sA
gL8QWyfDDnbx9ZdgwtcSoRTGkeSom+ucje+Pne/g5O/jrS2Rv4Y8O1PkrWpCDFqw3zOjGyP60HNg
VlWVwdynViyCuSzOq73TZ6IrCFXFmFDY+cG8vV5yXCzhfOR3neoI8zxQRWR8mtfCezDkqM7zds5a
n+76/BXjUAxnM11Ufi/NC+WVWhEDZg7BPs82Gm1pnW5gzAh5JnFO03lwSx1oltKAdPWUgXEt2BAp
Ua/35gDdXpGBRtSDN6nl8WxiigS2cY/nGz5JM9A9YPXuFryUGDg8GcaSx59KCruHLU7fh5Lrcxhz
e5+c6IR6PHR8ZzgkBkHmpHF2MbFj59s/1Xk4KRPm0cisVnMDgRZry41jRE9+p0BhUImKcVqprVsf
LTfmtMnw22ZKrE4TD2s4x1uJ5Qpg5cGGI7n+TCxLsaE2ljxQQYkbvJNRgEs7JsRoy9bzTNyHIFiQ
wexBFVYrQH7yqK72UL7ixxW2KaEXnyfsmAFFCjpZ7pMwPuFPvyGZ8Ntqn7i16LSDv2xkWcASzFNO
d87dz5f6mJN/KGUsv1VkBDuAR5JTW6LHqyz9e9fwAw6YNtZSmED90w3eoQtKzJqCzadOT5o9Yyo/
mnDWRARexBAnKWP2g7VejFHirYDCEGO08Ai3NGOz5PpMMwi7FAl8OVZmIe2mpwxUim2Ccj0gkv/v
ODeepnM3FZw+LWz8vXRebdWA142AJI+h5TUHa0cUYqaNdplXb85qf2ARpQ5ot3dv0rlb8kBqGyoM
XzNtuTZGCKmShhUg56mzK5QxsZ6yHcsQBH81AeXPb/vJptkWsYN8LubAGmD4v7eaKGME8sqEXcsk
Fan9ulLba9EYr4bkQ/Re7WoPODaAbw8LUVDVJn9qf1c+l7w5LjvVgNs/IZOr+/ojaP122+VwebGE
9cPKnJOY5u5zXsLKHomu0yBrLUkVhGLKN2m4oqCBjoT58QApae6BXB5+JrquVEhdYLPh3p+SS19g
em3anay3QdcjZan8ksHOlsdQwdh9CTaIXIPB5QW0NN13v9ngp1zkqGCPaBkJVRpFz1SsXK65ID7x
KZKgkENSVu3AUqkadmjbHHP5GZBTTdU2Dq0iala8dzVWmJM3BPG5kbHYCoFGVRDhXWK2+Z7MZ/Ku
DM9x5shT7k7NY7pZK59CHJmqEkLcyUcdEMc97mwWaG03Y8H6uVB5azqVHj4O065qS6HVmZgenKkI
UkTjERZEvGDdaPi9+JH+8hq1CDaRGu9GDQpTNe3DJQVlKGofIs1oCeeSRE4zpU1Xq2RwyBJkVbGn
EN6wrN32FPRWE89QAgh8GYEsGL0Ma0WfYCmFayPS38uhzVYcYAUXu6KSjsky7VyWT/ovMdkPAUh/
EDLHFnYMGjoGtMFqZCEf8VbZ/bsYQjvW3WMcm2aey1A4WkuuhDgMpk/gwRska8fnG+UsSZktHsBP
T6CwjI+p1z2EpTQUIIkpyjOR9wC36WzamwCKk3y3qWjuhPCBK0Yw8PpOZ4A4d7tNyI/0RxWZfDE8
8Yue19wFC8c3vydL6iAJYLi9trd0rkuokYfl2l+4BXZsyGDlbdm1HIqNJRGeY61WXbFlO8i0J96b
ogHC8l9IYM8VVd0irA4LMiauenHlbRx/QQ+OT5dtjI8SmGn30EVcv/fz6dStTytDK+Q4xp7Y7WT1
jwNSZpGuz2yypRRcYY6fYYNN1g+QgLTWVQX8eSVIl40DLSJM4auYGYF2dFj3ECY31bDC3dJgHWF0
PU5Gjooq3Z6gdi+DUfIhgpIOqh7fYulX9nHRwPlbzeDkkd6V04lffj7lsrQtVHsgG8/oA7xLeAkq
67Ua52Ln3TUFULewuDHLdMLSkAOWyQgzoKUZ6XmPsWcUDj+OLBHui8AgZzWwmvk46PIkYwLCD7LU
tURU/U4BFX9BurJr0w8/xdXV63xFyzOjtgBeUCzVk5FbbBX4XXz+/7fhyCrOk/iU5KKjEV+1HzDc
XwJfdMwcgnmmQl7Qfli8mP7oepaDBvTrF+xwZvAUFjxan/5uVUaZGIK4wc9mpAeEhgrl7q9P8Dxf
ekllsECNrd2X5lTILZnz6O+y32SVQMRPXSwT6OC4E9JPLM5GXCN52dBqIxfOcpsXMUOX81irsGtM
C5Azy2FrHZAxPEWR94vQE8eqximN2LrS0+fWBh8tG1uYGgnxgLwB7p15tpx893wWl2eGt2nskq51
oowkFX2OQKLOXidev2t+NWgwENHVD1i36CvGtVJmTNV5mOlVin9gQ7pJygDuaDJbkZCRdwwfcC2x
a00gWMLZZ2qWCF5KFb7MMybb95JwuQHEM0wK/3caMu8VLyyQaXBL4rP4luziL3JvT4qEteshE9Eo
aeg4O97zMDB3erVnGWxC8D1P3gyOcB5ZVMjCJDCxmV2JORZLqEjIZ37bBQUPrLoEZpspq+9aQGkb
kAevfsmwRAZ7LGDCTYTkf8nNrIYv34g0VbRONln7zvzARQW81DoPbHqhVX7ZSzWcbP+BiaYOtjrn
KRFIfL/hP1lD/L1fc79ZlOTuBVg2zmIL9AzCWyxlH1WyqdIloT+og3kQdcb0mjKljZfw+RVh9Vod
0fsYlZE7XfprkNSCmAR8dzyFZr0I3c4ba7IU7RiwqIK81pxGAfwsYb0hkn5TixDVVvoLRa2HMmfL
RuvhQpc21tHuWa5V3lwWF75j6rZ1JchRVXaV0dWU/G5U7rmWZ98gbQFeXZvmIq/0UVk+yXyOH78U
vIhvdJyJsVoIYakBSgWrEHNt0mDKe2oXPRBzfPgNo4/7NayC2X+Q9JwLicwBIcNlmvO+nhfvb34H
gFmhMs9LtykizPhPkUddCJVn9YV5CKSo+b7M/RA6l0NCmVREDTw9HDnRzrmpURalNLudO+2tkzz9
HCDB7+I7Trsg3w7ohCfKlzfUUQqjDISUvoQobKsYrwdKRzVIQcJUVrNd3taAch7rgA2qUJb+zh37
nWm+/KduUHED8kIcayEPOT7A3jyRzLXHeXLe3EKU8oxbF2TpVTaX+ZW7fpQ0nZnHkh6HauNO42ky
oEU1ZRkb1EgD5wQIg3UArPK8XDYcVdsyCE7XSr7pn5kjDOLlWGtXezfaTS8gjviIh7JURGA4P898
f9JdS0a6ewX1W6rQ2nn0Opf+tjcjoYLTXm8nxsdcxyijVyhSBo4AFOhjJQUR5xXpJsqmjnLMBodd
M0CHyupdrCDY1LYr5fQ3v78n5sh69D6F71UofomxpcUAr1RQJxfpF4T8pFExf1Ek7Dy0Ns4N6fog
dvcu8RRSJJGWjsGxwL4zKA/qECUPcrv2vmEtnFlAVK/Y76Zs4iI8zjcO7HW9onj/Ph3bmPXbnw7a
vXRf9KwrDDFklDZvrnOuFhdxkL7zpsq8pO7PPonx1Tz6Ri9+6sF9zdzB+wu8DJ9UJ1/MH8qinL+g
QEL8xBLsY8eOkZD+piH/LKIdXEP7YOwAOd1B08bvWYf0aeVp660MMx1KefhwaQ2m34JS9ddYj2G/
WNOI3QSazbJdIQS1lWri1HzL5NdDbZ8LWncZDZ02ywiU2Vy/5L+oJBN/P2xjdVw9avdnEHCoWKyH
vOl1F+WIsTUKCMP0alcx4IWKY1ze89XVu2ODMJ2MPr/PEgiOGkhjG4an6tdK0801/4w7a/aKOoIF
MPp/tnCOdWyFhqA7z4+73vLUawbZcd6T84y/uchxBxLA4dtUdWHp8KGZQpviHFQKZUqxoBuKkZJI
P0X9DbEOof3eY9jh3YwER+f0GGDkmIpLqUcwMoUE6TSiL7SqCZ/kDkvLLkwG1oVqmkVnPmMkfRcU
Hwyc92j085ekX83jJbY7CMAPbOEd5RHh29fFAZp2P8NVZJMd7rOz777uxajXdNf0JG60L0hlvBtM
pUcN+qc4Y6WA1HKkaJaOMQI+wB7+6W283QkxZFRZGFA2Az8c4fX1Qki5v+VWtq0l+Acybqa8zUOZ
PSq3xgHrE96jQtPXcV+IpYaQWpPGOPGGREk2MwoV6RpUC9ct81DwP73Yx5ueAPsfpomudeksi9vS
yCGDXKLdzTPWAT7V7VSCr6L7HCW2/y5hrP6uHzdh5QBVVJhKoTp+HX1zEhm8rdrbHNgnY96IlMdc
2pH9IdZ1K2M6wsAHd3znwvF5Ya7TSJP2+4uS3uEdhmzeEhYV1ypEme7U8bwqNy07F1iIgF0kjENJ
d9sfNZ+5ednhaf1XOa7Qfy2YnRHXBoVxCALnEfqGKl74Y/yeTR/qNFvdcJ/gPlnkz5drKaqH8Mwk
sGFE9JEqbHkTgUo7vhDLptpZRJ2JCpAXJUftsSSQgwmz895nyXVRkz9+/XhDNI3OQecwX5R9ecss
GVs3ukMDgOpOd38twOkaa7VLi4H2F9ZY1uEdkq86ULblUJJ4Bo6iSEAP9bizpuY0xkdM4gnxp8FF
+1Qqj2uoEGIPzcSmuqhUDmZ0wZvQuU0qsaymb+w571CzSZsHmFj5Z7tHivs+C7YCujdbxbnC6vdA
bQB9Knos7syF4b50C51nZFt2Yn0HqaeeyyxM4EAg69RAVkGPAztsOnVrbKai2C7bxDQJDDsOywyN
dKs3vgkqxblsC0naKgLLCdf6G4OpkEclF/1zfvZUV2BH5t4dm4DWttLoQbhBghwkmBBaapY00GaV
s/X+OnqULym7XnUBmNggXbNIJ9q6enuDz4ObbGN/LRbiY4cjojfJ0oaoqoq2gJYQ8GE2W8HCgGtG
kbTiWlUbdPcdKyeOtUsqy4ACHwijrG0C+6AdPSiVEH2NsC+beHNqsVEgbNfvvdQggAVuR7ab587k
73/o2sscAO3m6Vvo6rSWQ6/1Q/ScICmJDVbQzoC+jFVfE4UarmC0/drRAibAJR4IdoY3PqNF6VQh
fjGEzi/krSewHKKRt6L42LYuXY2pyoZIM1uSikNcLXrmLZ7mNCv36c8tKwbfio5GPsKXBL6/etjJ
G6OYlAKTqGrEKNgwrN9qxEG/jTp9baUP+T5TYBUOWO5mmxgkWWm2Ia3NfMSXJ3TtEQ8QzPbBD5qj
5klYZVZvDEfAO/xgtRdqzAIbiCqdrbnNozri9jUehP8Wxj0d/wfELfhoNjkVtYpq76Kuna0z+wYF
dqBEv9o8YAf16+qWLPO8GOvohRBOYhWvGyGevLp/PyexWpw7anGYpFbigZa/eD3fdEPbo5Bw6RNZ
f/MbciptGbtxlEPhNhfS8toOc+dwBPhDL7hDKS0ny0aEvhQ3PLEFfWICvqwQQaf0oyrhti2c3R1l
oobvOPSlrXqIQPy9k1dP5WsB6yM3s12iL3WUt6HnPUf8y9mFeL0bvpsvA3SY0mmmNOSOa/Zg1E5H
AsH5IeiioheTXzy4RzfgJlGT1RXdFABzyHuMyoDaypGWwWOcyw/BK3+/Gb/wlLPBDCPxu3ioo4GR
RNFgnmaxEKmaV9C7+bAKPud521zqff1KraF/npmhXSgoeVAJ410hcoJA51Qup6clwhjoJIqjICU2
mcq1i7pF92FQvjU2cXgiK4tXwFqBQQzxQ2ATQnvDG6AOIoDzn1DoftMbHjVhj1VebQOkKfKKr0Zo
mVIZ4GsJJk184qzThTp0cX6IUw3J+cYkTq20W0j8oQ9n6H3jcjxDa6NqxcFoAOW1IgnChUexdugx
JPo5D0MwRsE/wZ5ISqasLK1zJ81Ulyx0GKtiGo7KckAZb6rIjjVA/M/PoL1jxDgk9B7PWkT9yzvF
BZhsqbTGpWm6GKFy65dxGJV6U0swrG45idMCQBid7VyIxjMVIeGWFsMjT0mqvt+bo8U+CjK+qpgH
pyEifWlw9PvimGXZWz2//srdpdudifha8J5n1ymv/c2Sf5k0n+KIXk/kWV9f9xkew2wFKF+LHVWi
ZMCavhIUULW5kPyXRtMhWBe7eZDfwWFW3WJVj8ymKJzVCyyInQ3fpJ0m/FdL8K7YtLBc1p5rB29A
ioakpAMfv39aZf5LEoi+ZGj7nSD4YrzHmL4vdhg4Xmd8fkC5ADVXmN3tgELrQeRXTrnRH2NMeh0f
6PdlRMxHG9M2FRoQzMklNRU/AYvWOB9OTvrGt03P+XKqLxguwqh4wecsmDvV5rKZmyEslyLo4Pho
hHImBRvxG3eOdNozVw0I0fA9YDlKe2glinYOe+bNlNxDxhQRmFq6U76biZNzrI3wpOh+afp6+x6B
tr9xJpZA2ocgZSv1AeUdBMfYCqKciMQ8SayteFgCsDM0mAEg4vSw71n8C5e2fe2hh7PfIgjxlDgl
1A1A854ZV+k4BYYK/NMi46qXh3xLTfRLKaGFFCr7lmFvNTYirlswnFUX0Kc7VTlzY8pcyMVZpGGn
vjZPqA4EIAI+AOCiqTBsyJBS/M7UkXjucm2ZVmq/SLM+hwTUqkMRPe+84aXOybT00qs0t4eDYVHf
cdcPuw9nZuJ0dA8hDgo/2qLp2aUjS0kgfCtgp2klugGeG08vnV/NF5ixjy3BfVZQ81o+yW5euPtZ
zvUE2/rA6hyALRf2v7Qj1jKD+B9k7BGFI72HNgEAzzF29uOBu0PQZYXupOCAvm1Q5SO2AJXWHwd5
eHKLEDuI+UpWLwxG3aPjwoQZc+FhTriS6MuSELKtLtP8VVlVIU2Ld0TeG/weKXZWReChUq0XwsIl
qto6iwpT6oSX7Eh+uvILbC9r3HCRaE2nTwqQbavKHCb8bVupi438F89q7v09nvpDGNQ7rOPoIU1f
0DJhos8kOXx38joou7vNAXVGA+R8ZBBAeVyBpajIuwfiQCbW3cifmbsD91dzsnGi1PFNN3itvN4T
9l8culW/0eCmitO6gxzLKJuv/fSBzikjjkrFjkVdiDv8UT1oc6HoA1jVvT9ifxW3BklgmC/D4Zq/
vZtoWQcoyXZw93/JuGx1fgIOqZ6Qg6vPXdQcMCJUkBd22Dj0c0ciE+/7obRW4H0EFHUIpD4heh0c
AmqfCSM/O84ezTamb4PQHNbWiqiU/VPiuJLxmXzZ9XUhesfdVhvzTRAI224oBKMcSsDKmh0Jwtbl
ggIFwfCfejxPXohkVmozGbmPxpMcOq8SFYve+ffGK+i7nCrK+6swakXgSU6rIKwV1LxF5UUSBloz
rLSvF+0bFoqVilbmZ+vOXH5ysCgpPrdjhfOt/UmAjx7ZAup/qDFYJ0NTVB1vyPqRH4iQnuxH2G89
dp44DlMKzPpG5emLCJjPrHMfZwfiZXCJlAxdr/bpNc5s+P+cSqhcn7hrgFA0/2KZDpEbUEd7HSHf
IJ2pfR218F7FwClTrNeyrbI5C/wME4Gmxef3QOnRZVgCn25Jx/jDd1dClLK4fusat/H1UNay2a1e
2uLglfLtyYusW8IkUMvTXv7Yz+Aw2Qi5jmkOjGznAoN4yic2wgniY5IulhaJn9Q44mkcuokxhRm7
QkZCaSpWeTG6HUg/oVk/fZASh2ZgXllM0mtuliN9crLHfqN3PS/bNcVXc9rTR5TQEO2XPVqktX/r
uzxfW/mVTo3ZhPogWyvnpgFDrz/QpOHlOuXgMBRx/EONT0HF9G12EvbBLJplDyamDJt2cOGwI/rk
G8yh+AFwwZ/g7gmRzN5ecQ6/e6KzAe/XR7OycktwrBQq5B1VuS97iE5mV+0yNoATkVfhFWUIquYA
j+Oa+JBqMu2WeDxo0alJaeT/LzxbRGPWsQn+uT8g5jqlUJMJ4WntXPhvHDl2KOj3wJrIXmW5xzVN
RD+KbLsaofPcxkSgHZdC+6nUpSWJrFRPYh7v9hsnzolun7qsO0OyJOAPNltV1uPcY9t1WdQ+U6U/
t8wsW7t2aNaitdd1nTIuc5KrhZCwCHUnFFvFXpbIJKVuZ2pMO2CuG9GmfJ6xM6k4x+j8SL55PF3S
EmCiMHDQv0GRO25pGrPFeZRo1MuLJBaoP96TZH2Oa5ujc2ur8YG60IG+AoUuKvxUBqmUo3RgRuyP
+YIgTJ63DOuBFp37HkyR2gepWemPWbdsikLyiE7mb5TYi949gcWiFtjaHyn5IYgPsCoM/X725z9A
hiyY5arbG5z/m3EjHuup/oEY0SjKYPl5ARMqFjAy3vfowmPQPwEQf0Zo4gMUxNqxQ9nBZkoUdym4
yigV+eriHcJlG+2MerZlbRfbo81s2COUYqoH2shOgQhGirjssMk7vwc67GUyAFmvRqwgFxABjQ8X
KDOX//dvWMg8kws6DcmbNiGYHlGR6vf27+mc1rUaAY76H/gJVmJCEOKUJ+hBg+3wLyC8GJMPZm2t
mjp86vw+fACHvWPUtAYWpz/n2xrPZnC08ISNnd6KGFiT79hRNAn1BSZrpLWiWVOD4lTOAutsodeg
RVAu74xtKX4BinReyN+v2aMVyhSRbvgdVa9uldckFLl7HFCFtfxaBK3mBK7B/N4k4nA4scFbRFeV
HGb5f0N8s98RvjZFIWAxcEvJqzVDSRYXYyouSGtGDw/CxoxR56Q1EAHqSaKdqcdsSGm0R3QWyW+R
2mE0x+L7fa9L0sR9mTufoNV0zV0TdGjpFP78aYjS11DnrfV2RrPIo8YXa1Q1jx4524hfeymZWiit
A2d0EKhPkWosejcSlRNgqeRtRxD+cxCS3bAEYGGALcWdEYv+lJfvU8LDqdYSMRI9wKEFbMrfTDqL
6gyx++XfLXyYaWw75ntcHv9jBDGDFBRdETFLSONDxADJ27MB8Xas4GyLQJSMFHexNDdac7F1E+NK
c86gSOSY9Lnw9tBdyKXPTZ9Tl5yS8HaP1NAmNaZ3IKjIbJYrSKDJwHKsq5BgjFsc7AteAhj95Bcx
BKg/tkI5GaLTMt3sC7TM3TBs0alfULqG7JBo7c5uViKLVhanCDPkdST/ePG/fS2cIq1vEdVzEdfm
PhjSwyi6X83c9hnFzllNHJI87wwFoPfFXb7R2GhiyUEE0KnwaSwMNgJ8v90SJ7Fgv/bYHjuPpjGE
8cMmkwG2mzH0CJAh+GUjRv8lIsyVUAZp/9CP2OwETjY5jEh6qZkqqDdIQF4ctks4o05Q8aq85jJ1
Jm9x7N5pRvEZHnRre1DXEsOl4bZRzm5YPflom0VnvvK0sad5uuVN6EdrTvVzRdkLFp/vqffvGHd+
PrjfrsqyDKuUN+2tF/CQLevxVaDjaQ1MA1Z6pWX5IazGghSmfCRZ1XS+XWftvqKftnBkUrwsT6UD
afR7m7g/AnPJDbIA6Q/HO0ido5rLTS0AwY+AF/Ae8LgJuEVwWujpmFKuGRDmvGn6R7+VGeqXxJNd
diqkHIVAGvT3hThtpRjr7cHDK+N7mNYiQSyId1+6GfM7k8w3wp1MK9nM4LxkiBIX/BJpUgivwjbW
XnBRn84QsdeT3cexG9/ziIYneJo0ArUgqr4dnvNOD41SAIGRud9O8cLzQfofbTlSz+i9wIsSjGg5
lDzMdl6rjH1Vatx3UFoC4SQiU4E3q693HxGe3GP/bMgqQDqbo7AqwYKtmdzG9GOybPImOXCqqhV1
QEcBF+njIgKeJFjTGrQ+HwVFiknXMAik8FUAl6526+A4ZVrO+/RK2XsGsKlvPgnsUZu0PIg26i79
hYq76V/78Jzi+80lM0QLda1RkT5rO/ykjqhZrMUYMZama/rRUFhGSaFr2O0B8bIA9BpORTYI/GkF
2E47GgV6wBAmo33hKI5xTwcCd01xWSBqxIXPKxaCxTrmVP2/6zFZswUdGPzlUykUUXrmto7LVZ0j
a3Oni0/oRuw+3oKhMVtWd4KRkJX9vayDYkUaECjRk30Vgei2nWJxYJk9aG/sy6GV770f9mAeMdzL
28Xh6cipn3L89jKWnpecQ3HKCnwmYzPFvznqljT+jXHzLR/LKfE7PgLdk/LVT7AgzDToIc9cwc36
1yRfX4mtZPVHptYcpe3/xfBnO5OA/UjqGGCKWZYbm4H0qVwpuWiunihraFpyLf2+1ajBEYFRzkeO
wTCvf8MZQtrElXTBNkF0M5waVQ2m4OspfW1jPZ1P4ywn4g0VpcR8EgebzIKic8pvx6xikADGHtae
AHdo5Eds8WpQY7S0oSD4ARhkuMZjpDHJXdI0wRp0bzU2VVF2rwBsjl/JYowhAoGYvj1P5M5+cmIW
XASR+zXUZ7tpepS7CGm3ek4BIUoBvi5U/Z/IQUShyVS90oLbN3yj2gM6WAnKTz7iuONnKOw9j+TN
gG9qUi9D1gnXHwcpNYP+854ltxfFOrfRoHlTpVPEDXyul9PCm3D8SENScUnh+unuEhBRQdBBuark
6CkreIG9RXY3fY8Rr4z7s1OgY1A3vdGZlKzr6Py5v0N+5VjBYzo9yVxvhNIsY4rc5NQFTKLyHf2e
AuR6iVXPaGvwTZ0fDayOrmK4jHDlyMDd+CQ0hXBdiG1+sYLoEuGnNZi7G25pIv8wHJnCVZfj4y5g
ePBFvJn1rdOUAr3zCXkaH5VJkLbBnUvsHVhSXh0lXpqBeyCGAhPw9MpCMeDsUEaXvIARSxO4FGGV
4nBYT4pRww5bw4aCI+OEHpg6zn15De6zq1k0VG4eEXqud7PqOV7cVCSUxidlFFb86bUP52WdrQjZ
pbFQiTv0xSxUAZ0Xv1FWTe4QAtYKSDTdLXnmUx6GozPGYX156TI6NbKtGqVkY2wzHYmRmVE1cHc/
EG7W9osClXNX5vxnOZ6U7dOd0pKS9EDtvho+Ma3Q4qlehHXnqP/AwWuSrrKiIx9Q2/+WxDGiL110
ZPIbbh18/s7kNFtMGC6bbeVPcUBG2aE6ABpbSY3+syifZiHJ8F3zTR68ExXifJM4q1DkFZgpYrss
aCLGPEFOCyA3NhicqqXrvLEnb+vA+NDxGPnWiLaT8gBiRlpNWzW2uijRPHWsQBPD3zgDKY/ZStKh
AXhksFYrzSEcrxKTcSeviSY1zF5JE5Q4knSKz4Y9MBSG7LFafNIcuO/A6Nf/gkDEEbJpNuQkMrV9
L2xq9Jq63yV6adsbNoBX23/4CHBI3yrvcYIPI4EhAb1NvtmwxJCOe0N25XoftNmZ7hW/lmlouGdg
ijlUymyzCCvz3TQbxpB4hj/wIbJsw95fhU6rAuixamXPO0Un6UT7GDNEdwPPaL4WqqAGukeKMn65
B4PykoGYfqcC2yc8dprC/oi2WMpR81EcMoMumIEbhJ9/iIJ+6Swq6pe81t1fzIqrkWi9goK0Icaq
Uym9weTbVD/HxvCvkncle7CO3MXeb0waIFR/wnBK/YZP92GVP2qNXkpVwrleCASRQNXetJFLxQiL
2U4VN6dgX0wMlkxnvWZqLqtvcPg5KyJvctnn/Z8M9xn38hUgtq6EvxQEO/Mc1fgOJucwf+7oAFww
b0M5VNBfIS9wZXLX5aQ3xMkRmP7otD+9zzGTZy1Qr/i4A0S4oQNyoQvICQIh/849CDF4LzmO2XK+
BgjBYo5f2uujtHM9dOB2tR3HB1tzdn01vSyMcEK79OsiMSn4+1HbKyHRlGOtwGeu1RAB7HmjfOpO
COQ5rvMKUBZ6QxPrz1qihmCV5nLf2iNv9eniON5rZnmOGtan5fTiU2pmAsBqU7QWf+7gQG3iYwek
tbF1eq1KnC3X2yrXmTspY4eZJXj62TizqWcn+sGrcYP8uVHNuk4ndwlY9KxrqTASEOlBb9pXh7OE
dLbeWRQUQUzFY6f7zUyNYJ5vHsZtoEkRQ+cBsMHe5prz6/OQYi8zXWCqxX9Vby5qT4OssZnyvpPS
mSbTQida0kZ0XDWmASDB4U04EOZZgn3Ngrbw/6VsjBS2Id0Ez8YLv9ojc0MMmQaGH3r/wC/WrD4X
kr7ifkvR6C64a8G2lKq9ccRQSzu3x8X8clBv3YEJTZMqcvy7G8VICiheQ2daeio/Yk4mgGfVX7Xb
wFoaWsZK6o8va7DIMGJxZP1YFf3Tt6GkLEjmu2Rn3VsjX/SmDcdfR/Qhf9jlYo5pQyn4vPdg4HW8
+o7b4MeH08W/ELqKS2YKPlcLeWtV7oI+22sAY+L19FgUIB6KZexrioh+l8pQ0RCfl2abYMdSK8tE
BkvGHpAs596mrUDq6gm7dhNnZLtC93UNBiNp+zM9VYBO/2TLjpBtK9e7hZRVXvC75XN/cqTVDyb+
p3AOh4O6mItB6f0PRdPJxOg+IY89uo7NrF0RCu+3HoGqXnDq/hFIcIbb1REIqrhEIGy9ITYbZQqR
87Ed1tUFbBmoLIGt4p05/wsPTCTgMzM49CeOLGCPVD241qFaN9zZuASy/XJCd5Ur9MTA6Xq4k23Z
s1dCKuxmUClFtynTLM4bJjgeTIEUL0VSnPHena+Cynjv7HJMagOXPZG+6mB4iGWkiFFdUP0WLb83
S8va88VOyF7Xf3IXSiKVh96Sequxf8Ee6KxPvHSUsetfnQ6ULhyxte4qjYaCri+c9gmEYumBhEmW
OLCWhal4WS2GoNtGIBCMPH4hrJr3PIMkDHPmm2ly6OcjLnDuiDmQgqwEM/xF4mTftkQc1gtWxhga
UDfs70hO1gm5upAqb2UFb2S+uHzx9rGkyOp+oZc8R2ROc5iMn92sYVfr0aSS7ryfLk0WPCI2PuCP
fsVMTYCh9GCv+yH0yxSDysU9FC2xGybiiD7KqLyvDE6m+O1iaZ6AvhR1LTPgfS4bcacx+kvZSqHV
5XpUh0U2KHNM/7wU5L8/hhwDkL+BiuX2BH+Aes6JsmZVLFTEBR+oYlZlqVoJHDJ17LUE/ToGnGwB
KB4tlftJoWNGvPG8JQHpVIoWzm2xLHuIrczV2E4bPy1IGjkzZ4o4Gpp41Z8ZnqkdLJpOkyqf9de8
I25DDq7fgc/KGKnsZXT9okkIhlGvi4FAjlCCjjw/0Li2XimpUzTPvuWBbVvWe+6DEALyeHZbgdOA
nQIbqjsSaAFt43YABcBUPZjPEHrQUyfVil1tML1dEdbU+3ekCUFqkDyjAAZVWyNIZ3GzESSSbzZ1
9ffQ7QLrN3n3uSHa9V+J7chbtB0fxouHSF9I3QB+BF8z6HGNUKE1kXUqBH+G3VYssogF+bRWzRza
XYU0VYGk1QLQuX+V4LNQaAUv0JCmc9b6IokWTe0xxKH6gpNfGuJmd/BGb0czHTdgxPCaSUaW1PAY
72NRV2KxY62HH0MUHSk6c611qFmzT4duXdP7oe8lPkg9z/ixJydO1fDkxUoy5ntiUyeEKA8d55Yz
1YL/+dlXRW+a2vLlFdprOv6dIkF9nVJHcFtqRiGph9MYRpor3nPPJ++6m81Z1AxT1+RfhhDOdIMl
DW9FbUB5gAyqijvIDqQwJBcACudkCATdkVAoDYLZ2PPiRrRQF7bt1U7ki+XCg3MLO8zbNPwQHjKo
f6O4eHYhn0pgaE1x5T1xkywH6UdLJI2UQvCUigDZARLwqOiSYl9E86WX7A5FwnAsuWLl82AgEp37
PVruw5O1f/ElCAe61eNmL+aVX6gpIC1ixbwayM43ti/NkG6VPWZ5LrpQgug/YgFeA+4/51xJ+DBc
lJOQo31BJ9YoGr7hGzisoNiE7tybIjaRABKNUq7btYrIeyeQ3s4QqKEcgpcC8cqaoQ6O58kQIIp7
+L5iDxgkOeYfkN5sgxD0bPxRuDZCW1NQCNEPN8s76BfMJjIcAf933AvcGE/dggBHVtw08M2Sz+pT
XSs9uOjFMEFVUP+Ri/OUB5MfLa56486+BMohguV82fJ5Zx60MD5cKm8o7QcnYW5v9ft3sNDvBxp6
7xwmGAYQlGm5twgmShJnharnj220j5zt7L6yeiNvo/jLifQ0KVPFkUK6g86JyHYFaI+h3cJ+snQA
HWX8b+Y3tP7R26Hd/hYmJ9c72jxAM6juCpsFnUi+A2y4uGbsS92d856kpE033qFJLI1dHqxOFeSz
ZgIAFRivSrFSqRgtNxPrE2hfQo6vmUQ3/MyfpDS88tdaYSfdB9Ig/maWkZ2yZg7xnQ5Tjj3hi+lP
lIMOkTbUHpdkbUGSiQFRZgx8x1HatgKSPbjol0VmE/qmlgvAFQB8Iwct1WB64EcOpw24NKMawZvi
PuFHhqH4ymTWXDfjuimKgjgqbFrWW5T8TpjVkecdIa8RImoF2ui/6/52M/q4UkiRZScgXzbRm0jC
5hOvZ/jQ83zYDC35qzZnbu2w6tigxtmnPtAovIdRWomlzLfwSkXKRQT5H9NltyW6OPXPvyw5+GGy
ptONC/m7tCTXZZ5DKwLpxwqLi2Qfl0uP7Lb2wKYOIDuUjHofgq/c8Vs+29hRxSfJFFNHtYBH1PO8
kEX5VCMetqTTCQUp6wG+aRiwuIMBz+cczJgHrtdJ9d7oBtehbwc4Q06QV/WaXXWTB41inC7zs8Zb
gZP2kaWlNlT0lgUvmo6nGoJLLeuXZbWgknWJNxbsMPB34WmFz47hxbNYcW7riwR7nd26z9kkbJtR
EPR8ExVTo5dlouSqYbRINAQOLFneO7bVoi+Rss3MZkK6PbV4/P+L4YonamMYlfJ6HrpsMRAzzfmG
KxVTKlNarAc2mhlSOQG41cigIlyi8Y3GH7y6vcZluPDat1npIz/2e9A2/dTuR/1cVC+GPYazLahH
TuXeUbIqO6n6UqBWSb3XfUMzFFYjO0VjInEgkvyv3HhYvESMJ9BX6JRfVhCk55e1c+sIm29CJDr6
FMCiB39vTZU8vVXmpvB+MsA1uibmmIcfL/c8tX7TUidouExIOQq1nrIRsOLjBpmAdPXtuwu0U8ri
U/TXvAY+bWCJFO5t+59Q7Bc54ZUf0STdZ3PXN9d6c3i4bomxYVWmlJpLl8qkB5k6XX0Xd76nl9/K
ZArDJZxIGNRMyNIOdo45ycW4u28QxL3JmSxkhpfuOS2g5SPIRXn1PM4qf6AHY5LcyZcEfudun+Hu
FD83tSC+MPOqS3BYrqPPSTMy1cByCq6tQvmwKcr4La8owK0DfdOP+JDNnIe2No68LLMxq1RLeon8
27BDTul84b4FMOB3vve7ihGU07Uz6CTPDqCix2CdQetdd4zN5fJfLvtguFEqYI5Wufbir79JwRT3
U5tQaWkWG9y9Y6tv/4f2Nt6XGresnBd4wWCAztV7JoFi2j62Ct54/lMvstKZqq969tJykLjqeru+
EJrIypwnnqRqThfRZOGXOzGix02DbnWgZ5BK3FfXYvzeNchH5JKI9P1N2BuZiDIH0AZk5SjLxJAa
W26IrGZ8O5HZT144SiJJRbN/ty/lHnfFyywGJtmbYa2p2aDuKs9VBLoVgj89LlPFy1at97CNLRdn
puV59bet7YbYLE5aDAzTZCzIV9nu/SOJIwFHoBs3Iq3A46Q/rOOAj6xoBXFHrP/bFAxJt3iUdwRD
R3mU+tossfYM2VMkHBu5vi03evP4bQQ6HI6JIq2mp3VVOVDnHawl7W/TXgLLHfK9+FpQVvGZAMUE
BjEWuz8ZdwoN6BcIa1QqMJg+9iPWzmu2TRsDBow/0SDlVoFJ1CjWw2ysLF4fnqHKjKc/vIrzCtcN
D07TNhJ8t4FL4nfVGgv0q0NgtLv7u25LQuUNw0M5H7+62aT9Joel5J0EzQJLpBLlyu52LtEFiFlW
j053EHhMsPT9+ConKHxQXhha4mzGiN2b3SVI1ku67+orXT294ElcdxyacGIxVdPId+h0iwuGzO2o
r6XQBucnnKQx4vWXyRij7/lRTx2e9q3vQBTzU4eDMVUH0o4IdC2vMSYkkVizk3bL9mH5EYi+Nas5
gSYqQxjuOEXS3HRo6M879QiEdbcgYk9VwVlb+aI3vwgpB/qz36xqh8Q0EGUv0f8POEB2oDaIsJde
W9frNqjfKTBlrrHbH772kjGoOIHy+xCZLH7dyz8wZ9hEvEg7uCqbcUiTceUVbgS8WaAp1IilCVct
GO2bbo7sz1yYacW/KkgY9ehziON8wEujnzIKEzH/I1vCYfQbB105vx9xiO8Hy1qQlQG+YvC8k3Jq
WGzVNBmHOnalv6GBBfpzyHZdpYUmTT1XLJ3IJuNL4ntrVzmnbXBHESqMfG+wPIAIad/+/Dg/UxjX
kg4GIfwUgtJqUSX5qZCqCeaFpYy+kDj6ls/0mCIa8VTSVutD6AcMZliCw6xv1KIY2lzsUp9kLDd+
+Mp60FjBhmhNAfUnT0vAiSUyGGrVoylLiAjW4xperVyOQUww0cTwa+uvU1Jl9UIRXlq85Ed8xn0n
xjmTlBhx/F//4PQyLAd14dxq6ELLSpg/NtFRR/fwRP7Jt7djbBvOaJytKJwq2BpNn4dir4ZeC2e5
Nyyv5yGm7PhU4cUkn8NdjF+W1vG+DwgiQOrPUjm1KD2M57MnXJD4m8rd+canNDA8GShN/GAihVft
LEuKbft+74NlL6Ugbv8iT04JY1hjJ+L4YJMOwWIWgGSBr25za+a5l9mb6YtXR9ZfdTCjDP2Qzf/c
PuNLNK8mYhMhQWpUmOZZFq/e8bTDmAsRscmuIAHBF5GzsTntFXcuhwz+xb1Z+Y2fJcsfllzXrOGf
Hkz3D85qc0CkiC5klVuFR4lbhtJ3TN+g6IUZhxg7H6rajPB27u2eAYrH1sAovXVf6PoLOtvRdyRg
NKFs9qBoJtjyfjVGs2MiJnSgtxQ2g7+PZ7q0hYscguSdHoDhL9YC7vt5RNTANS3i3TVxTy7qn4kp
TGNEHPFGO7hHIUtCTw4le2b416POHI73yDe+WJgG+5RvMR8u2bbTCyh7LhP6KacHaJVNBfQwT6z3
5YZtTpX72GmeXnSj+ZLkHNtnrVc9kS06i55EkAeNXG0yNs+owqOyAOOVKRrvIQhjtZVzB13L9h0K
sdDQiWYj7Pb/pOvb/rwbPppmrE1p3C8ykaXMVwBXAvMDAmIGdDGysRuSm56xWWY58IKMNBuyymMp
74lEkP/w9XbU7N9y/h6R520G3AOoqEPeEH2yYRGJNR6wFtY4QEVDNSmOKjYxKvEy4hFz6VmKhlOE
FUmAh4Mhq9IFOhMq8fFEDz/3rWnNPwDuLtnX9Z1WGM93kk9F3fh4LYTiijJgl47sO93/cnl/xL52
lE+/tGRD90pZqGGcZeoWhGcoT2kAgEBmUk5PIynClbtL4IhlsAtcniGVh9TAHFITwsywjc8IIGom
X1WHSoqwXIf3GcMLR+xSBRvT4JCYztgc5EORtsuoqO9msyIGoix5dsjw4v/0w/1Ci1/tAmR4Mky6
Xy6rljy503S2QLIuFyiXU3MAduClFoNwGucGCDdsSWmF7j90AXwMs2y880NId5mZjP0IhIokmjxe
Q/8G2+plBnEO7wolJvPNjVADrfPW5LjBkJQo46KncmuyOv2Khj3RlHwl+Jmxtrslt4hgfbxkvP/0
9//5PPWqruEiwgfkBY3p0x9cTNrIJh2uOUN13tBTOc/8fOwyotguJx5BKqfVFjMi2wWdG+oaKx4d
7fw1+jnDkjb+xKnEY4g6YZTTPu6zlPaHw/Ld18lvnNlGD20IMTemQFoeYjyo7XEE6RfFaxJUN0dD
0n15zP5LNg5NyVLnSSBsRWJw7fs60MRVVkTJZV6id4PizWcJWQnO0BgnFYivpIC+UfKnVz2gOXiH
/IZga93sVwpdLKNnqeTIsHqWHAAVosrrfMbrFT29Q3Spbu8WUxTki2bLMEvVSNmC6JE8kbOarDBP
NBgQJJfr3oVtbZRN6SdEE3mv1BsI1byJu+VPqijhxGCOpwRTmRUeRHMMRv6j07V1SZQTpK+z76/8
M11ljHJIkD6f8xp8JKbz2Xzi98yvKuHJ6BfGKfpLBOOsVPegWsk5US4tZ5NpnxUxgSJpMg8AcnhP
Fbc0MqfoY7Wen2dRwkc3P17wFhbhh4Q/JKZMG9hOkhsQfoKW+Nt2opyop354Gw2KuADCWKodjtCq
4jCZgbVjlUrH3L8TReYZ+L/K0Y3NiAk0DkjlTuqDo0ZMihZCgCs9RqY2syuMMjGfoQw6iDtlpKK/
cl8957tt4w2XMIKoF2+oWfCy2c+2tPb9Lb7kLywWyBomOvF8dBl3tEIshR5iZO7sQ2pdONjJFEZ7
UXdP+dTmZhjJBhh+wHUk8UWzdB8Fi8pZH6vRFte/9RHXeObDY7gJGPk86vrTcArt8N4OJxCE4IjX
iQolesrL20g72emeANnkq+zmSh1WLIJgNDOskj8/YVJWYOdQ1JFtsGutXMyLJu6gHpOTlI/00I/k
3qV9DNyFVGLKQuS8LITxPm5jWK/PVaVEkhv17fYQPraI/VbLcCEtzPP88Lm0HrTHUuk3mPZiANvK
DrBvZU/LhPhxvZXGlr8e4EHMRxDyyiH2YWvKsz2VI4VQ5QtkaAfHwY61Rkb9Yz4iEfCAY8Bkt7Q1
4dS/JGeuqRp5uoxu+S8Jrkjyx54hhpuD7lOe9jzDjHKGOKUMa/QR0DYtZF/adTTgZ7YBVnbAvHY1
AXUOUM2iHF5vE+uZef90asDhnijOay3Dtgz1jjUP1/xYkvR0WtGimCgPfPODu6sS57yyc4fgfrKT
5e1IS0VwlKJ+OEp3GxoVcgLuc6Urt6a2wSRXHWlAMUIssY8Q3UP4PgLMFH/hoIdvQis//8i77pXM
WV90IbOxQY1ZMlIpCl7F7D6dQiIUy00Jwq/maRfpbPSmTZFu68TO2EjbraCPaOZ6wCS89RvUBdNB
GulMzSFGgyNw1Nqfb7AHwI23KH1jPApF1IwTNQT+La+IxC2zt45rooF7XsQP6H5yTHqzcgyFEEIH
3fWcm1BmHAApkdp2wp/Vt4m8UU5xeX3jIlFBGEUxnibahpQC+1S+qRvepP9svZyuHyVb7XT1Tefq
5FnzQ1vJph8KdB1CAn7XIaqWNEqlc1ibDlZOogPDiYApw6zZytvbKFuW0EXyl2m3T/rTpCzrGQYa
68c/WeVx9wfn7BnB9wcMJ71rNR3vQ2WlTZlMftO7lkc6dxiojXVUu6E9x1rXGyu+/JVf3E24RgKu
gnCSdsfgsx3orCJDxnHt8OPrKQBsYQuWXJPktNuT1DHvrbsf0JAxQCJemfTzhA2eQkx0Rik6Ugvv
1ixvB9v/4n4bmLxCEGRfWe/Am/8wdaTm65k4OsTmyy7MmJ5CaYOLk8WVZ4cYFpJblRvzcbZBD6sj
fPewU07PB3FZrg4zxTAqeSbK6+m1C7kKX33/vFd4QYhdgdAjjO2nCew267b75asVkUNCHbTeIQDd
Nfh7VjpRDt+GAIiCWc8cV4TJcxmGN9vU5tSDJg50GOay0b7c0VqQg7lN2YGwyZYkcMdtVaOt9thI
Rqk67V3AlDftaTjQQneQ9xsvSa1gkJ6yS4jEsnH9dDVG2hEV99xUP1P5RiFVSfV4ILWaolG07VIE
Pa8CaJtyyHaaXNAjQGWklKCeim+YpBxyciIJ1BAwYsHKQI168j8chtSCzSh2dvg8yOBQjmMcyJJn
xYRVj41W6PM9LLgz7KR2oYgZgcBY1TreMYv954D/3dO2oAvRjirv1LEie9Y3Y/GHrBECdXiEReY3
6M0HjXpvEhqJrBpV256WW581AjssgJk8ZA8aSykDhCwH7Fb+C9gUbb4MbfcI4h3KbrKfYCxMDtTO
rjb+y4T9vQ9qWul4hLdsCMJkQFV735iEgOWv5lxgcA1h6SxVQtQthyfhW7+fsvci+xPQPGzlMiUU
N254Ktn8+zEC8/x9S28cU7ZQrzbw73ozQkxHJG8XZ5vn4CditIVLnXkdKh5OzcyHyjZiyJ+JkL6A
MuBZ6i4vxMZGBfOAMo1EWEmR2kHION0n/PVjCPh+shdZXr+TQYSAFT3N4zjXBTlw1KrCcdIWWPkR
bsH+QMHlaRk2aE9kjJYPrKXFrgFUyBlPEOghggrR25GTjWEwLNg0R+6C303ss2fVS5muHKXQ2AGl
TZarIx1UhHJ8fR2rtIoD2waLTU+j5N4onwgeCXRCF/GsJ8EsGX3URoQqQU3kD7AkZkniSEIF8gP2
qyEVYzmXBTlfnm477AgTzFqPj7WcA2jQpMfViYczQLQ5lXo2kqXoAjq86NkbqWRHMW9NXuPaioCk
fxSU6hku/6jW6sfeEf9hmAmba37ZCs8uF6GDmkptGgxE7NtmUE8jfzcw94SmQMws/hGEgHHfg9gY
bluUIZfBH5dnQu3bcdlZq30IwonthMaUq7QW9P7htWA+71MhPrpDSvujbTQuKXUy5fOfqnKSVvEv
DkNQlhTiVVqBeVCAwNdwVl+ShHLPnUFFxbqzb0SuCTBIrU/fFYQ+iWPiapv5f2cMicIxNXHzUkAU
ZWaQoJX9j/aL7xYpXFSdJj4LSX/9Vv3BzYp0T9bhqmnMMdIiLHf5YPEASIn8IFJvifIFWtvHp09f
x+3tcJwcrwckI5QpseqllyaII54sm6OSdYwSPNqDWcPUMEwaP3fryONS0hMAQntQJZAtQfJFScUt
YtIhQ6BffUSO6qqqBZ5MqDT2E9H5gqyr7HtPF5Cro/FJKj++NwwfQiD8ukZdbRHH4AEpWT/v8TUi
6f9y4xYdA6yMjwPtkQdIalst5Fitrtb5ypfwMdklN3JoQ4MOd0Ni9LUZoRL6S3bUbmre1TA4J5+a
r7xaeFtswW7kxTWNUIjwf9XqwKGym2ajp5no8BfpGlwGi/4gSe40+wBp4Uf5GE/3ZZqJRNeEGnb9
+L+Cr5U5n04mMPa8yx9gGYKYX0sGONHEjpzObqf9+z7GNoUfMehItrMRhXwoujcvvixwMGDSN+CY
k+GuJsITWzcmRuW9nJ8E7N9jVhNjlWtWmkdQdujmrC5lln5/W6a6Zv9qFTEE2phQNC+HJosEcL8i
FBmkl/GFoSny9QP1DYyA6q7sWEf68atykwAElEJPADLJYL8AjZHla1obBBz8w599+Kmm1RjUmPV4
weNX8FLx56qd400xS1Pb+GzOzLyVcICd284XNfumjEUyWb0QZhdCyMWYPquiaDF4AcYwBnVC5e9u
qqQVEDsehMBW2FeuBlJBLIAWOraHVHRRsOVz10Ctydwv7ue+yqg9g52M5Q0bWkMKRs/TpEbEZN9d
MSlXsxOLK0d7xFwSqbw2pnekz9IZPZ0u1JtW7XR+RjKJ8Y9khY867V78pHd74rjS1h0AVpFdUV5g
S5tFgKABTeBEgpSsUVYlfyv/0Eu4gJ1+SVuybHJq3cswWu3PVVbSi7KPAsFAXZwnNhOq5rRmiMeJ
xQWK7hZWAlGrnAXqOde83nZPxNGW7quYBwwFq6OrbYnTh6ERwR6qmIWS4rsExfZJ421EZT85R21v
cqNlOmIFrP0NNzGXp523eQuoxKEOD6UpwrHxmIRoqufYi5CKLex4DNBkz5QxSbd8EDNn73zMVRU+
lnW1FmguzhLHPSy8ZAF0ykP4i64pQd+F3kAQvb3+YXhtwjJbgTHg8Sq3AFWQ25d3QrBs4kSvLiKo
mQueChYZ9WTy9NwjdBDmUOYuyA7zQs2CsZtmeKHj7QtOXXxyi/WCY05Nd+/KjAa+GvZH8wjqPGrN
wlguABv3vJTJ0+MGyUg82F1lXgJ0pklxSHFkTig7EP2nEnCfHMMDQfuYkawgXkFb4nYvDVTRQ84W
RMF5oDW5j9Iu2auGjLUX/P+MIbZo7BV8yH+7OTV8AUeV07BlCWy2zQsSKqJ7o0OSDSqVthdkJ7e0
h9xTHK6siWmvx1nvIW+97sF7J8pEEuDusmZkrZ/Sg/U7JfTLwIjqGrMdL79l5LH2gfHNTHqhN0Q2
Kh8W4k4mKg5ZVnPC+5wkhXkmLS/aYa4YosQRwlsx5ZCo72pn6woRJfCdIYl1ovOXCq21wKKB3Gj2
2Q3RclpbgCoUnG2V0Y9GwiY5YtWb7nZRqelzQiVXjheOP0lqZi8WdXSwaYLKA73DhBobgRS4J3UN
ChDTVI63ZT/7SuQvbv+5A1gqziIGi6Hp7WkUoWzKnYt88X2Fxov27YafWKBddW/FAKXrcPpCbIYM
vjFKBZqYyqVkZB9I+iqCbnxkZ8EJ4JHqnJ/rVqdTCxZoBjKY2UFKvSAKtMPczvmwnNhj4jYrZK2B
AYLkdEfav7jnz00oqrCAPnHcIrvtrmU5WCNmJMu4gHXV9D0Kal7uo/pkdiGARqbTDP6f4NNHhL8W
Hh7qqMnlEeNlHyGiXKHplQacVJPTV1KBX23wZkRyEWWPUX9AHdJJYjz30JR1EeqWT9Ly+CIKz5iw
dokZBsX+3ZtVnoT1Ua7Yco5XWQ+DPCY/DInOayayd3ugGhW5+das0ZpCxsWHsS7r3HXLDnnmV5w/
QWtnL134PC15DtXEIGRRBdXkb2kz/1uP40wx2pAmzsjrDI7m+ZcKuAt+CCR+FLmJfr05oVksyO7H
cC212Yhi0GuFspXv10HYyNCSuKpS14xEMZzTAJrPg3Fr+JrHZw6cz2bidEDu0VntufSkM41krkKn
pjUMVENF48Kfk/aF+0IEu/GWijs2otueeEnDDWVbrypMMPpKScZ6Pq9OCsJf2+hXyXuI7vMNbnfl
A0aa1JEF4u1xolwy8WnsoQ5L2jdL5ymyP2x1hnMEi5Cs4QweJM9sZgabsLf5c/g0tEjkN2v3FoMM
y5AuMP74otDIiFyRlc/6yKbCXElL9+v2+NoPNEMRSIYWf+gHxhCqfNxQHFNGPvu1DqEdxO8jZ1Lx
5l8aKkC3LAeVj2+M7PHgQP31wAD8Q9P3dvq/n9o6fPWdhQixq2JNmJKOnhsUkOg9MTguRHO9YzPk
85YR9ioagG4iZOrhCFKG5azE5mctfBV1Kt1DiZE6fAhYU3Xn/iFDPdNy5GaH7/Jyoacky5dJXfvG
S1f3wvImhz2chJszsellJBnqjr/ilvyEpGyP4BcF6RbUI2Epjk9ANHAfiCNPPE/WxLY7MvEsDrRy
n3gIA7DViJ9nbQYoVukeoxQ48knS7P/6X5zDncQ7rmbN79vwnW6+jmK6i52MgEqhxrlnV7MvpQfp
p2oV/22RfIojUd4xvfwT/MZniVPMUhn052LEls9gZ3RmlC66btzHAflVqEhGjv6WBIQPVfIWGz9/
VaxrqmkrEzvSRIhV40CvKVa1CrtQmhU6X+dspuLJtLF5b4yPIg2i8FvNuLO+P9bUi9YrnE5Gzp3o
Eqo7m22laFRXY8AXE0yr3DPDpNOXeT8y2ygIrRCz8tNsiEJ2gUM83vQk2nfB7B33dhXNPiopr6Ud
taTt7Z74f75yRPYksFJi/dEc6IoBpOQksLlC4HDXRFa1d42OXvqZz1L8gVG9ed7E2raRFDIR2VHx
Hz+K6GzE2XREuwPzqpMwHvh/YcpZomoNwvSl9VTusM78rij4WvCJnA9T0k035Mm3abwmxBypt0kL
T8+pVxOz8Bcmve6JUoGU4V/0OU0aYIsw1eoum13UIe3v7nTVuyGup2d1RFP22tK0hNhI9kgJXHtk
HOsK45yeE6u614lA++JJfq65/l9OA73yTOUN266nUfW1WuFd0Jriut7g/6g0Ox2yx+OWVquApFdl
r3c4drTjPEBUWbKSX+8GI/GsQGTQZKYZEY4DN6kuyIYB4RtTXPylb7ZKAcPwcvzBG5OVa8+WQOtg
8w/PsrtJhoMROKJUmkRnbwrKB/BdBQUizZLtnGdHdm6TUbxsYNUBs/5QBcm8/VCxNIAcAQJeouaN
hwtKcSfS1206FtJrmrGq4QepnWd1xZZqWJhYBbmuq9x8OFL2Trm5D2J3VSyJM0xk0//36jYKEV8j
Pwe/Hg5/PpF3iXEXdR0dM1REBf4rrDcz2e9lGkeUW1RGIwGc5VBVG/nTTEjORma01pZ7GIPinUyu
5u3nUN575iIiRBwQW1dxOW8J/OpK7UQER1YKUcI+fzBc5RRHwtJtya/7WM9crIK5a/i+PpYB1nib
JQmks/EWdBvINmbxq5zrlhDqHP+JCgGm1WNNTANyIBCFldqHyS/3Wg8d4XMG0Y2BSsIFkQVrdnI7
AXHwJr+NHAN72oMabzV4eJemgdsODCIbe6kMxwHtZOjac7zDTRYXqTzGiia1W1uvNxL3bkFprubK
Pg1DUqyPi5QnNZzKLfFj/OjOJttVCP8FjAcNvlTaXvv5RfDPMSz65/1oYMTEJdEKYlPtzTAxueGe
1DDWPY5Y66dEOCgJ5lb7cW7XHP1fKb2wgNFSAm99SBAS3QcWUJ3gMK+vxLPwR//WLegHwASBi2EV
5Q/YaL8pCNvyTvqK76H4oTnNtzU8mW2GDIX2/LQwThByjGSyesRqweRhg2auEORxTai7MG2/VfM5
uckzIunAapdtKNMQ1fXkSYO++TpUzbBabtUNrzlr4rVPRauqzfnyIWmC8peopHmgjVp8rVByCYv2
A17/PneeV0IAh9lTIyeTJmUp0Kj/w/2BCUDA0vPr7lGTAJR6/b6SlSME+TKXZB0U5pDw+KQjr3M0
qkOwLxEwYyU8lQzIQEGWwNcqCPNWe0HvoCE1Am4GM6kbgNS+V8gsNN3qmcMIi0Cdtao4vL0pj/B/
sfpYaqQT659kTkpGFzrS5dCG5d8ynQi7Rjy2aPGxtZJi5pa9dvC03LyOVqJqxM3Iw6Z/zjxydh3z
F1GIn32FB5sYalWx7hqRtf9gkhlc4qTKiRhbTH1ONF12dxj4PEdl19SiOkPCI5lEXVvbwym72Heo
rYkBhGT7QJTASExTLxztd/UNHq9+uxhvlQmZow4THMDx39bHplTSrluAy2PZsH0Si5XnF8mKwGEO
Fkm2TVc9hkt3r6dhXNldUEw2AFRT0bSAPQhpzx5hksaLPw5Y7qMGN3LeKzUMJvbqOzdgxtV6NL73
GXt7UWPRHIzl31O9lfx4eFMLQSuoMtq97zGio7ZKAm86OQO8t2xWC9UR2wpU3JsL3osZa33hTbzp
/eDsOJ+M5VXg3Pg6gVyrkZNnuyRzUzrH7mdZfxhyiZLO3J1JBz2cgtnXc5SU48OBp4s4Vm2/PeHs
EEX/qe5tSfQ35uuMWMQQcvSPfwWhJ0VwGYeo/y7VI/Ds7A/eujf49VHienzLiWRVGridrGFp0CSR
8ILwvXVvpxBmWMPME9IzOM+d1ydDay8/1jY8X8wh4j4TS8Axyolj5NosTYC68f+yclgh9vLnmSN2
tswhQHDfCDA/sLvRgPPKGMh/Lc5lJ59WI1DS+HSKqd9f1weqXu/xGC+ZwS0q0kWGRWPqFK5GqcLC
brBCbtrgYBo0sdZ4+SUiMYYxIE4mKL69fs4YCBeHkmsE/S73vYXEG9zXOmqXanx1eSqgdhq05UUb
Yv8p6ra0xMY0zrTYIOha7B2b+KEzlqW8INwhf4+tq7/09ujiTgOR2XA/WRfErzNGe0FPLdk69IcU
FnJNstuTRzZ6mfH+qqX/+DfqpjqwqjDDZs4AsmHdvgpthh6rRfMkKGfX4+KkWL+cc6OFV97ScwCV
XgeQxSyc3LetQ8tXj6MrqoEfkJbSUKsOl7YT49v/vtvax7z+rwII/B6TQOFc/oKJa6OEznBYmaOE
M0KQPyNeMyXYt6gCgylUkLYNbRCqEz4aUhXCfKgO42WJ3hwHBP1MSX/Xty4DGK+HVponR59MEz9E
YV32ycwEY6kJU1sD/s4/2td5vtd1rxTOOPZHQyj5uiVrCFw/PkJ4oIdUvA07DcD16ZNmhPDVn5W2
TTns96c6L6DYhFNjwMPpmCUQrg8Bm14mwIAFuGp6pO55nloYM5ZQUGJi+dTGsXVZorkA8IodQ6bs
kJVU9CfDxWyibLNRRlOKHs/oVtnV6nxW2TDd2cZ5NC9k3y924fS4hQR1X1neJwt3WrQKwRTITheW
u1jP4X4KRiDtWzo9O1V1mYGKccd5hlTI1MVOi9fWrUMakES4Lzn37lFntaClISzvPWBaoo4ijODN
uZq2KWrWBFkVYgj0/miLyThLwUNO6h5SL+t9xDNb3ii+8FLOtuuN/HNBrnMyhJ5P7w53Sy11qXQ3
gtjXc6UTNUMI3QrqptTv2gIxUXy7I2O5nhJtr4Rh2D+2K0/fGe4BpgXmJ0Ok7tVBSJx70MXNZJe2
vDXeOf6mG2Dmcef6ORLGm0Rtg9m2LoPCVdahB4H9C+l/IlPaslRr46KcwvgbH4nN9uWddgi+khnE
gUMsaRF6SddIsm+Nze0Mng+7OnkVFNxp6NNntsigtWZ9Ct8XzS8SmUWKyhWDrhugv83zV5jkFrlD
gdMAYDTFWD5pa1OGpB5gbaFjEwkt0I4Q829UuYoFvlBCcsSkP9OKvhHPPT22HM4/5cW7TqrMB8wC
4T6nP3lsQMo9aDwSoq36i3+h7YHxwGPAIX8DPAW18D5GViVJFdNmyTNd6CCBlmXs+uJbQ0qZTKjZ
UvwOToIbWfoIYf+kiRM6+DllGAHNJ/CX0dDwoTw17Nwav4+gm4WfGmbzk+YSpzZZo2TRR7AEMpRC
27ICTzdZP9LN1042t40gbYUJ1QiA+KhzXhqdTLP0EJGmGCoiwNwVUS8E69KMNZznoGdFkqk7p8+5
nDv9IKnvT1RisFyV3w/MQOFZ5eFCbNJUyZ67+FXE3R/kVTeuheG2KOXQPcl7SXV8Dx75HV8gnn57
0O/WkaWHSz3cM9Fnv1fCmGDWgxlqZi/VHlRXela0BRrStMCsgrzQea1vw+qzt+K/7rwAaMSs8/aT
PNofQB1tkVy8OvU6D5RJl0NyPAdtnBwhcb2K1mwluNIi+jo6nULQ+KYeTLQ3VX3rQCio8dx+Ntyq
scjM8wPTrNNaQvSmqmDD0goi6oHNQo/1+/Cad1B7K+/b94K0YLOLTYd+pBMbics/XeAAdwhjOUrR
hhwVT9+id9kotM3FCD5FV3LZlk5ZtKUht+ypximKl7lEJSDp/W1EfpGTdUzBs/8UhvhXdHbzBCnB
7KQtbMm3wTsxXurlT9Td37vZ8rRvwDuPyVNY6ps7AwaknkNSpcjECMJ72HlSC+NRK+SCy71uExMh
GA+MlxrneG8BRK8Iz68dkH2LrVP6X6YqD26X71laPGwgiN3sDbLvUA1Z5KvtLzqeKlRW6czXmniI
e7nveIScH+reQiySvw8e5zf8UVV+IpxNfDc4dBzZAs4z2cjXqeQi4Uf78NRcQxBfIEoEJFv15gom
89gLnPZId9gkO9gmOYtTXHIcAwrg2+T0uZdl29fOfohaj4qIEPRqBGuhlMJhJR0r1VSCPlp5D3HO
YzUGr087bGHM6sNtP6TMoBftViAJTQcKzQzBB0tVv9zcL2T3ocDfXYAQV7C6toMpD0yBNSNZqjcn
qULHolKT6dbvCVsiM8lTLoxT2T1xLnHYSNLuQYg0OAA0Mgfp66gk7DJhu60ns4coLtBfkBPYPkP2
vgheZ4zntHbsG7FxKCMLAMm0S29RwI5H46/answTv6nUXz3KFofnAxxC6UfeO+Y+Yu51w1ihG5gl
5GUaT1D8pc9BBYQKMwGF0xRd22cFrXWF1LKIh2sAv1l15wrBw1bK6mG1bhQyLUNogLQMzjh3Q8ES
w7NSBEFtZVgBar2aFiVY9MC+f0Vdfip3zB8lKjYIaC90ys216/Vey6S6XFpIzDw1pHc4LD715jh1
057MTSAnN4Vu62+GOZCPfA4OBK33s6lZuDgdj5BA2btYRHb/bayaL1WeAdRG3WzbrK9k+wve8cua
BzhdoL7cKDX1hpZNwAnqX2A9ebIEB5bUvnDANMRKdQD4VO8E6q7rFMLYHmmZZYoYU4Q4Srz4Vv06
8RA44wrAxKR8mM4XYhA4yljaG4wOGw9YuMgwBJFDqOxn0UWmxSRjl8TSyod+Tf1af96ipoY+ywjo
ZjelArjuBzKrnyq5QQuOJmUiFuDY60dTZumYdFyKHjL/GhI/ljZxc+j2XdI42gErV/9cqD3ErSXM
fY2HhAngI3GWuidisCeaxf7vtpRW3jxH+qpC812uBFMtWe+wkCI92y6GOeD20c0lXQ0PN0DhAjlU
x2iTR2Qmasu6jZ1xh5ztkXeBJwh52g7dWK/BOCeYFLm8RmLW4JrHW1UuZ8H4ZeE5lPCFoPvB0knS
kbbQnUbpEOK5kgw2mxOQA/yFej6savrdUYOHjpoTQa1xEcSTlo/4m2aHiZ+Z9mJV6dBaIq2sMYkz
8vc244TYmUeDAfzccYTRk+aApfDBvXWmvKjz0Wb2hPOcsbRgKArBUqdfZlmAqEf375AxuIjKJ1+G
XjjlRjqROlfKKsdOeH9z5/2qUsDZ2jpqrVgy6SkBYNgV+C/K3SEDrSwTBhLDjwfmfjAmA7XsC9y2
Xmh/eVlc7G3sZOktdmWJ9vPOU9OQ6hF35dTIpfIiLh/yNXG7O8nT8go/1SnMHuX89et5PMrFYc3o
tF9Fqzzyvbu904WeAzbQp8DQbCImIuXjATlPH8ifZvNbTzG8kdggVKQCCCXtIy8cPschregPJYXq
PAWteXS9QXSQQm/7Eif5hhndPtgC/t16mEvK6di2UzeVu40GzOrNLNl/NC8eKtOOHSYAbGXtI4y4
eYfLJ5eW28vA0rww1UHqD+W0YjV6GLEg5j92Z14/JqifdCIZR3QKoQJLIj5EWyobTMi/JNeGTxe9
SuOrEzB3vXtQ9qLydNGk7w3p7wjwjGXNs2M/jfcF9/FtwAjYQFzotCjHqz8vv+YYvYPQiCQPz1Ls
BgYz92vVuXZvR9XDy5uSQtETdYqwGUkt0H/XuvKYyckqo1N/aTX1j71BRwukH2XytmjHGKg88Sb/
FpH7MSbIe5QCQNGBpqNgGxBS7//ZsjH2M5wW3yj7jbFlcaEeZIi1fkfzWwfUT6Lq+Ewaik5rJjll
5EsSlhGm4bNKdaBo8zJcZ+6kxpqsKJTUQ7Gcgf00DOofkovm5fExkNOkmgfWDaqV53OyzywCUJxW
HG3ENgxGUzILgV60xfa7fG7vDJbgG8oSQSiMH2jg2qct0tPOLfaefYJzYUL7tsRdL0tNaqrU9mX1
5vg3arw9NkiRDC245aZvzEeqQ/mO0o/MuvWYKn/KE0CeDSIKJWE3ljGRyv9SDOEpwGu5IPuJbzQ/
xJut+nnQsxVj1EAhWFQkhGPBmnGgSGUnyKfJkx1Pmh2iNpvfVMzpNhct9hQ5atk3sNu+GKhy+vTg
5ys28ZzTIIGbi1CZRQXJ63VD0rlQynyRaRmXhykpJzYmHhd61E4y9OWtDP3m7ldx0AIfdNhs0Qqh
iIOVPI6FjsNBWrFQ0Wk+6U+eL0xQ+ajNY40CAbFaNfjy7abNdGwibe/4l0MMpNs3aSyDK/JR6lQK
pNYZjkubK17eLC5c7um8P2SesvnMjK/B0h3HKDFxQsFq9QRNf+j30HG7802Cn/+JHjtUYNpX0IJN
+8cVL1gYxWCEtLwKmRbOP1P8ebyl9F5np9oMVrDte5vefbDbhTrA2Hb71R+pP/o1AEtMmZDEdYiC
J+FMFNBIb3bEj+4hjhCv9o1leIsVo/pgDugjUKlSw/TrPcEzNpP6xjGjBWaVeKCHJTHJ8T79AjcO
4F1iTcPT/HOoBUGmm6nBCXgzmNGTrCuDRkOEHZPNZmX81O2Gn3r4QE/Cm+iMVBkSQJgEvbFpo2ji
2JKKJVJgpXNmltZ+ysXFGcdyFFSVXQKzbO6TddLOPqiN3CPV8Ksgan0q4FWcji3et1rcmhouJid1
FdVlT4cWegOTxiiWwZa7kKNw54zuWb5iwU6MQzFmotnyW9hrOMTHJcxJBhKbPIgqdlOxWGuCzIKS
QRCdD4cqN/19zOuoK9rDG8vUY+Xj2J26JdjkoUibWTOaUACHz5noVX+09gkPyoNJhtUUfHcGn0bw
MH5HXnD1BJGuLTanVJYsWoxerQq3O+8wj7s+3HByk6gvLJklIS93G7201XGqzolgcrw4bJOjAwQW
JRxCw7gxWdfwDLlC44MokEXzHF+LBMyc32ITYN40IJs7lNyHB20mRQzIZqkhg8xMSgtgu0Bz7xp6
3gVcOaxKZPA4hkUXt0JE0kYEol2mWZAYbOOclAN2RD+aEJeipBxDD2raMSZMEAEPgXjxxpPbtG5a
SKOjJMYvuulQbhP9UOuIqhJ9SwAe8KFJSdNawz0OF9j/D0t16OI8aPMjDpo6+mr5Ji1FsDuMqJEk
daQqlc5QqzPhzfYsO2QbK+jq0YY2c5BJ8BkqySLP/lokmBHGu2gxHZLfEOGkoInWDzKWc7zdaP+f
LeGdPo+ulIDvy33s4ns1Iisw/Yf2VRWaSQC3FInAnHk8aQLFAnAQZzzUV3hWmcXn7FWTDg/yGOnk
uaZ5VnUkj9k4JEUgkpBDFb3SKiY8I/RHcZUVllt+kPZbJWUL0HRWj/fI/WFOF4a54safF1PhoHd9
NhPDkHzcQ9pLCpjmfaO6jdq6Ldj7xXvL/z6GpiKBffYiA3tRwcwGqCa9iqxOZlbfyNGkCSi3QuUA
RC1b7F40hyONTIMCum/dGTKPDdYEK0d08QFv6CCORofP8kzBVcD6IzEUqOzWIDBlhmxSRukel/P+
pLdh+jAhr+ypz9AsxIZEpM19lxx/q4T6AhZx8/5r1b+pzw3MliuTrWkXPuZd1yxlXSs+4wbbwSZI
b0pwELd7mgLl1EtxdwRdVO6geCRgUXW8zBTiHZPilT7SAsc0/yYFFPKJ00P3mAsq51Jt0KCBRm1T
2iffRd7fidQL29e2QmYH2pLYESv3uWwD8xk9om/YbfODJWgr31XfZzB7PbjxKv7EYQ7wIH6LfVm3
l50/D9pm/OnTLDzrRcW8lIxWHJ8qZU6eNlAKnDIjuqFquvEVwe6jBuDDWAybVlaStefx8VLiT9C7
BCF3JsU5yO7oxCYeBUbDV/RVQQnkWR/DXl0vWnB4epEqvP1yMst5KSULOwBRvrCROj0UjtDSt9ZF
R+u4k0vh6G6qHbHWK29vJqagh/Y4DrwKpcka+kMEd9z9UZ6yuc9TxQ13r7uOVXAg3SeEN74qCLkF
HRkfVUwRFW1rBsQyQZy375xaDgXvzFnO7OXGhyl/KaDWb7pmlNC99JrIyMpI9hzCJqe/xVhphxUH
Au3FqzQDi1WBhdmJMj1pthSozZPn46uoWGpRLiiehp+TsUkOvaOrjfyX55rrtIQzlBXSMfauU5hF
azT1niHIyWAMyNfDww1FxitlExZeTTPHzoL9/eNeKcL8R23MBrM6kdC/vad+upyb5GA6nKaffZG4
6RtljtHTJHUU5ozo2MvQinzbeiU6FjH4GAHMHsbtHGA1IGtHntSNO7VSGJQvYW3F2DNSGOipdWJN
DEHlctQDcceBsbdwkMaagL4uRcuqzb6ykBTPsks07cf9Hxc9TCBTxIHY5wUZ6DAN1zWz4vvKXQAS
BHhFvZ4wvY+nG+rF1Otsyjna2SmG0GNvgRX+4XBrUE8o2i2acicbaR4QrZxn3ZoP2CgenPs/vUQD
LcDaqNaOpIsX3fcuwY79Kb3uo7UpdAFdX/3+okgJbdwSzb1s1AXC+PtGZZ+WFYK1SxKhn349qLQ4
Z1SKydMvwj3lMXn+fRk4+lRC/nBqaVwVKMhxFG/QLjZ57LecTkzZ97KlNY9enfm36iyRlMhtGNCc
ysXNyNwHljaIPJkLxffcaTQv1v5fypkGp5JVZBUSQW/PgV4ehRxGj7zJY7JNcQVg1NXApM2FdBJi
tvGpasy8Y3pPZbxLGPt/yZkw7ohAdDd+qUXv/fvg9vdl44aZLTVdy6lH18Ydq3gxHn+T/aOysWBo
8Yyfp9oO0EA9+fN5tO71LZ9un4lq6ozxwF/qQuYgRjwzY5Pu9jp+A+3EU9XHBPT+O6tWCYAO7eih
vz676FPBy8BaSN5Riz9qeleqn1JghnFjpwOv3CgkOXMUTfv7mKIta3VzdjTi+7Z/82vG+vhoidQl
kbi155Y8sBWogyGPKvrwCTzveXOC+X83Q3Vsk5edEt1TfiR8ZFvzPwXLWwPa5HV8DnCiQcMgqGjg
gXJ/H+7LLzg59rNlqdBni9AVcQwZXvpUVWab2AUfv3H0Y/sN53emHWvOoWvbzhqaKOxgQRfBQp5y
xkCYmvmJWpwau6BNA890SBB0eZElGxVSW9wyLIhwa0E6xki0swri12b1IPORiRe9kG1gMNaM+eLH
1apltN1LNUvW1VviS4c+8TVMx9H11BSAOXExkjVX/rhhlMly/17gNlObM4maAZlBdzH7BsBpocmO
LyB1IACz0P8SpooFpEQo4BrvnG3BDa7dEZdHDc1oEgQ6NxYmK7oXY3qMsVBYz5mnDOaVWzRvFPtw
oRpM8DwsCmSWDNhNYeH3N0uscLTqHtrr0nV6UMmQX/iVLkbkAk3CMa+wiKSf+2xScHSDf22QJKVH
gwYxuj3YzDz0bLM4/sOEkLTpijVKecKPKxc/ckpUI6mFI53qZaK/0SNVDNLaPdl9TD7pNZbXx7+y
B6QljA7JmuOx6mzsRYMXXH7Li+r969aat8ZsOZ205aRimIdzrvhzkBNAfOHhCIgjtcpz5KgBL2xt
L/ZeVzrSvQxxqcIATlKSHQm9AH/0MSTnuUw9lJQ1tD7i8YA/K6Bz9qJmcuTFfbOVJRywddZGl0IA
SH8z0BpL+GrILVogb3f5b0I36bvd+Vd+eq5SxGt+k6gb80lkj79aRUuNo2ODkOujkR2PnF6dGq30
Xivgf+cLl8arLmuNr9oKC7Zz2uUd6EZzSjIxgnLPUAMAPL7w9SZSjmDIZ0aPlC51eR/FKkk7DQJ3
S1QybIIs+ymm5Ot3j2DsTcr7SaqkkZ7Emx/Wdv+9Rga55zK+lDM98a/3hUfutVQB41dgvm4vUXaN
/j1z++7xY4fYODnNFaEIUDa4rRiuGpgJKrAfP0IMq6h6lnWP6Ob2Eio/wnE4bNtmR1U4Bb8GcyQ5
W7JYrdjl+2nqu6GgtRb3zMgBtDtwhbG3K4J4oi4U7GT7vBmciXoJhyx8PVYRPIqfYYwtienPkTtq
qGvDqm64KnrWidkbvevAIl+nLr2tg0x49p6syVApPJHrzfHJcljS0k2iHggLPCBeeMVdlfh4oR3r
XxIRhw9fQv0J1Uh14btbGvSj9q6jSpb2rnlFzFmRoqZj663CWx/PpT3ogX8Z3NRMkFeeJmF6iTM+
6jgUcVieWuph5Nc+9/+tQGiJEUZD/MAXAI0SrVQp2HtVakDzC5tviy3utGkRkfaZpXE32e0yhmZT
rzP1X4Xo6Bk5daQkgaYeIqrSKSRYmwbwoVr6HnkZpO0OvswyObormp5dWQaszJMu0XDkTyYvmD7A
3pkzrNE6vyQpyNSbGEfjL12LHZ/mQWs22N8csIWDsaKdXRMXWA0ti0FCoMj5Q9Fq4xP/XoXHAEEQ
070K9JUNWVpQ1JCTeRGMPRvqkWsZqlkZiCblUpKu7iYYyKiudk4em8Btn5YhbiuEM2huAke088DH
mIpGoVaPW80Pxw3i2GGKD+tO3jSjO17paU1tZEx4WU3qB4T2TcyR5d8yxhp8ZjfI3TrQgTfqImE3
0g3WZ2uhLxhhG5x3Ggjtod1FOT35cWy0ydCfzWu3uB95DGd+iU7zIlAtY4h+KIezq/VhwWMaESYc
D281Avlu1dGJOMRkuSQZq3xHdeUhGLY0F5HiMvl4jg2xq3DTwWUl4tVMtaoPgPtHgZh9pxBiOgN4
8bZUZeTHBoo8H3VvNpL+gEEZX/Y5sAO0sSoD41sboMrdFL0W178V4CQG4zqO+8xHzZrIvrFaRj1k
xFyDRVKnIs+kWMN4ibGz7TXnSd5v2Pmx8PfQ0qF6EEFX/Orh+k0CDFW28i6Xl1BW7EiZsxCc38Lb
9ueBXn42t/xcQYInnilw8m72mb5kZbBSTGZfVEegWHMD95BZlWQlN4h0e65hdB2rdjv1q6yADwCR
wrScIO+31jy1jveoM4Buw82oJdStq1TbayQnr8aAbivEgJi26ifuuzh3LlyJVx71K8BPIK98ZQ9B
0zIdzUKEQJsTmqz8tBhkGok7tV9lJntC74szFE5EooE/CEZPUHAsE8b+AD68CeOIUuIHmKmEP6Cb
S1x1AE/4bWvOoabFbOuE8P4EV04uSfrZS7H+/o+lWzNYTx1Zc5jkjlPKqtTqoefSLDD2N3TyotIJ
RYPmAAJyN/Of8byCH9AE8g4i9M5lzQJykM8lnBICaXhCau2khFmjiK8cdSVEVDj3HNGxFnCh0xM9
j5ojJoNRiUrlpR2M1esny532zflbIoB55bK87wn2ALm1IEMZX91GGzX5G9DBoan+mjnbX4QMkexp
Di4jo0DBBe+M3a2peQbeojSiQBLUuWbRnoq0SltG4Aa9PPzHN+PBmon7I8HUQjln9kXTPsF9pBNM
o2c7bVnZlU8FvZsxnOOc2XvstAgxHc+s7IYuq3ut/bB9Roo9z+wigvp43XYMZn90jHqkcwdmCUBB
GYSmYskVhxbyezQWcrL8X/mpCD0OZbvT1dZLfzA70oNytksiNXdt3a5Kb8a4nrnz7ng66pjJCtlp
JKmEUcTwqhAjDYIZIs5PMh8L+21vs28o6kR+jlWrCjOfauuFEIQ/Jy2nxvP6/yOInwyNplV/kdhQ
Z1zHjxBSHUPPY2cQUfuq59dQstq3KqGlrwSYTWNtx1WQP2d2hbp4ZVmrAMoZVWQxhJut3pE7nMg7
IN3UGmn3BQLkH3LSy9z8hE4TsLp6suUl65w5fwkvDJAGBygRZH5//zHm/U/qArIKFCYcutVDYRUO
IGusfNmpC0t3k4NrYg10/VB5UEigftFirqmqCGdUjMan/YznDnjnqUg+6Q+TIWuLrPzO7wbJW9Ce
UcvTCfqmbHwKwo/Lfq0HKrSg4ms0Hb7mJXCmt5kQDD3aZ1v9J1rPJHMrL288GRncVMDiYysUD9zO
Su5UrvoTRDRXVqU294+uqrvtH37Og6QW2jnfzCNfNYEuSaWO5FxD6BV0N6i0elQZvrxh+CB0RNkV
y1ki+OtauayTVVaYZQEOno9zuIi6mUMSgFe4IjctlNpjILoYBFG7qhib0y8W5Yi8apitkJSjQaiP
fFR/JIS8/BZ3gzimMZVHuQRcZt5+OdeDJRXHSF+6nHJGXji2aZKsZw/d6BFqI57bRTGz/iQ3vK3a
zjwGHNLA99LFu9ZDWMtEZtD6B1rWp7prEmjgu0rh+W0I5HoY6mNATwWkCnKxGyeEsnt8vdYbf8p8
+D20BX5G4ROIGW9HXmEqZavDvNQo4oHnUCbqdmGDu4l3XKgaYGJBemAkA+Vo6uee4EKd+nOkMLEx
pazILL2LfeL8l03EYTjB9YMUXBfSM/oFy5/MoSMCkc+2zRGR36nYP9I1aA1xzhMLzN7iPNbEAPUV
EeTGqj0w5jyJ1fCKUC0WOWe0N+c+0BDCyBcfKyFbqgsGl3Knl0vXs1I1FbW/5/LOT8ErOP7TrwhF
GB5CzOOFsgrCGSBHyZUsT33kRo/EFej+zMSw6STSsXfNf1qO6SQ69L291xLuDmxRM2dNpZaTUy1A
mHaoTDZrmqNfqShu/uOr/ycBmHGrUCLl0M2gE8/qdVwHb37k82fVHJAoMpebErJ69Vt8TA8j5Pfl
LZbkO5pfWbhyi2I8pZt7Q+y2Bb12A/MZxZvnu/jlduJSFSUfSvEzv7xrTzG52G65fKQLn42dcM+Z
2KAO+dImazh0+KQ0a3FJDZmlRNfJTsY3c2BayucOplG5XX15fOvfe6tQPHikafw7YgKWelfl5tXx
CBE/aQAmwibCosplphWiPcSjLgWpatWN8rG91ivYY6LDRUQVSntKpvFNVmYAsxLUIMFrI5TqXSVE
9+ma2jRnw53a2tKLrlDi3W4d2Jm/2Cebu7iVqT0YIadTqtmz68iKnjmgqjVGCuilFMsXVLAYADWx
QY0ODfWvKhSvKg6NZ0POQ4F3ue1jNvYy8VwBBlHkdLd0BotLs6nBf7NwxOs1Sij9Rv1G0rfjpKW3
mBNIdIDo2shWFDVBtOL0S/l/aXo0w/k0ubss4G5lW8dgnUkXEKPRutsgLV1aIxBn0LD6r0yhb17a
//JqFhdr2CDbhZMD0UBbuACPkAzN2c7iq8UmgLut6DVA4BqjHvxu+i1hCgdA/FnbRSNtY4BZDDk3
/E8ioqABQzNnL1pdseGLgUm5Kaib8jCVumj1dDG5LYKgT9Fn8ZlVM6kwu+E/sXSuwD8OUXCxMlVb
3DilhMfffO4UhZgr5p+0GrgkMuMudAIg/KJNRnCnuCbuZj5HXUwOHQGYzhz3MxHgvZMDKMStjfyc
yc8Xb8cGWsoGP52A3rEU+bJkYT1K5NeMBWmH8OL9WWDVQmgpcUFpYeSY6gj0YsGRvb+vJvdgZlZ6
udpFitShY9xs6TLNrC/fh3OeozbS7Q4GvvSknTSy6vpcJr0alB0gCuF4ET+/X9iXG/oEsLqNFNn0
T9iLowhijNybwWNEnKxDwOfqxEWG5LlVxS+OrDUuZJSzpioe4Qru11LKpqfyPLWeU24sgmZWqbGS
Sy1pqgQnMHA5c9ZekmPATt5g27FUt7+t1pqw4T9yLQ0iczVdMYfq9ubO9BLF3QqRUecza03Acbbe
M6A+FK4vKdSk/2f2a02i5IHoXHJGREPeqLLYUu13ZojOFa9Kwahg9LsKzowB3CMugt2VwdVrbVot
BvVxKwzh1+MCpdB0z8blQ/gKVkQm1TsvLevKpmKkfuMrUhNFep3qvJZ8AYD1Ss8kiElcWihZH/Au
69b9RguitQZtWPAfdv5a9UjzBPeDq3U7K4upEHt9Ra6looqsAaROAyApGiQbmFTBdUDLz0bxdBrD
3ZXs2DCyBoANMrR6suBfHwxS+rQu8bPEcXkGEw3oLuD6x3QHNA2+M0hhyaWSW57scj4ghqM/Sjue
RqjzQSJgxBXdjUXdZ+fW3bpr/sawpC2nNduYOm7owfLOY9qYtbgfto+Fuy5Hx3XLiMjuUpgKLzcN
ls6ESv3uWMhwiC6vJYYrFWh8j+b3J8Rqhj0MTWoV5BI5GAG8PKh+zF+BmNkz6e7LqRxHNsEdWmZa
hmI75+gZ/7BboRtX7CM45wstZTv0kpDVQoG7N6tJ9wNENotZ2z0SHz0H1btlny+XZbEcG7EBru22
cXpfTaT921EsU0TWLze9dwP7bLEoJxUmCh97v5xDJcL5Dfwx1M5SH0kdgHVOT0+Oz0JSCGGlDEA8
pf6N2COJffRTELeRRXAXbOqp9SyADOiqS6kGHzzlbrvJ4X19TxLFTtHRrCEPKzHZL6Wi10WlDYTF
mC+xGJ0LI0+LQRuZNrtc0wVmJ1uIVjP1CvBvn93QZpZc2s88LTzi4XcC07tbOuzqYGZMk7iHBMuT
HjLYC1Ga5RD8iD0wYG8P1oQ3QSapkux2485f/DOH3G8wyoV4Gh2ghD8dT4ed7wuBaMsprnlF0RVy
RHGNWohOKoephLcWBK88AhbF8GH5WoK+YQDGdYnhb5g+JYUGQP9k+76Yy9yVS9YFpB5+LJN0mSEu
8lVMzKCAYAt2c51/Fg83J2Wlsk1FkMTNi9Hv1lrfI989opLs+5WsL2n/YeLfEJC48Pcu/zT8G514
F1xq1M5s1ZM3bec+m3CrU9S1aNGNA8hq8sPC1Rq3scwxFqx67fzp1uf8d8qPCB//sOKrmB6e74ik
3z/zP4cUM3I7xSNM8SPvoMor2yy6IcJlxa329B1dpzOHjtuvq0dEr1fDdZRQKJbhA8lTF3McpkXk
ZZ0soi6J6O69ODKqreQSvnY70LyjwiX+SrkCHrdVvviT00QB2X0aJDSJHX5TNomU3RRF2ZZlJNG6
skhX5C2iVycnx45WeqzHtX7BkytXR7WCRNeK4VsskaAcouW6HByPDIpDdB2vpbgq8LP1klR1DUmp
c4couKMSDc6kJnQRmQEGfDjWjSWipDqXNnCei1qVYedfUmtrDI/dFupj+oR+8bkRY/bAsh71DMFZ
HOiBEX5XmLtvzrYbAJjp9tp93QuP7/5L8pUUnZxGiu2zcshMX6ZYbXMjZU3B+hGBlHhpJDjN0i//
+vYXyZA4zAZWTM4hKNjEOQtFyD/KJXrn0jVcoJNnib1XvvQEON8/OhOo932q7pCp3qy433bvmDPT
LJ8pUMj6SWg09yNpm5ak6qDRJYZa+v9ug07LewddS0WXMeycS+10ZsWGUaVZjGlXtiV2jIAfKRhn
Jn5NjAth2huU5Nzfs1ze/utvTPoWuqnY7oKVJ3xuwIjm+XuAOJprkGMBTqnoJPdYmudka4y41e4M
hQcVChJ9TkbM5scoN1MTI6WVJrV5kBOZxK/IArOLsvwkVpVZ9akzcVVgabPlEs5BVrElMO/8TFt0
SYhT9Qo30qwuYRU2EXw2BnwJuR6jeLZIvVl1n3H0NnofyPrtHcHZoJP6cFeB3X3Z+M5/2HSyBUQB
yRJVjifIvs7mgZZ6vGSaE0A3c0NCeb7hroutZUnrfgtiGJkNVLs6F5mrAC+gsp4T9EYk3QyzpKN1
l2qN4IzkzB4p8JckvJ96/ql/kvKb+o+GuhillrlbmDzGRHek7sQuFGQucPUBoyYBVawCRObXR8OT
P2Uxe0RXjwrWBY8jjMAzlUS3l84sBrEbM0dapswBDOQp5e73lfRpbm4xc/4Dc+jwB2xGHH8lLHGZ
e0w9jJwTw0QT8MFYeRtZB/0eEj4GHkT/G6XcaJEjo8Kb3q7V0I4VqAauywm3nLiDGUuuM5egf11S
C89stG8+KGOuTdnIy1UlWOguqWoQD2qGUxkTP+RGBTh7eREZzqwxyolqvKHmZRK//ZKQNEEZYnTS
wHOznImb4bwWelr4PXwZLsZ5OdaFzPNSV/Pl7ZwZub8a3FoNCtNWWTS+4fM34d7SoHXdfNH1kMep
3AFpv6q5ctBiZ4VbNOxhBe/ERRJGmVn4gDkd2fXRHBsNgnClicgUkjzupGkN2dHgrUVBuFWbVaq2
g56PSGRN1erjua461dJt0KN1LlXrmAQVpxR5SP9xxk874i29sbbv/U+/AswpuIP6XG6PET0NwewG
Uvxb6h+6H3GBuYZXje3GfLznMQgue69mWKD0qsZiB/hu/tJD6YHPxOtiZCn0kHzRGktB2Jzwd+zo
PBq7SIaQToE2qF6idFK5esad+AEYWLkwfnZY+DzTpxVeNGMYK0fTrhN8G02NPICCsjgqF/fVDaFf
vkyMCeJDQnq10vbfWZ33G2hW5eb9cotB2onwHGkg3DLl2Dk2WV9ptH4KeTcuB4Rd94Ufuy3v6Ra9
hfB5Fvu5KXPHEt3g71RLULqYyNVrFh5tEPMoCXmKKeLAG1eOfHY5kP7njcIg/QhKx0Kb8G+rlfIs
BGZctP32SajPdH7/+5eumJPjrwTu0DniEoSKGcwJjIcpQ/YaSV/PqcXSa2dF6pCg+ypIoFGrQ5Yq
jEMW/j648Md17LvKtO/AgTVMU31GQoYyPo0IBAYtD4Yb+hP8QvkmdcV23n1m7pmYpen6DY6spu9z
63/jnE6rWQdmivvbx5mKxy8BJoeKfqm7YeIXvjbhCX7zP7PNFGuiyO390io8NtYG8Nmjs7KW4rCG
Lmiy5PBXpOqSj5VtedMDtHoxbEeNp+w+PdZCbWMkr1Dkl/euH2GkQ4z4Y7cpKEpi/4ZuYVZy42rq
W9aFG+SU36vyDq69wXDcxmqBi2c8gIe2vgZBFiZqgzUvpTxcXlRdZYUfddePYqI96gFsTVKGxYCK
/hTmC91eAakpG+zpLGQQsozDkiL4yBbulJn8Q8Rge7NLOdXvAScZbFsmImB+rZT0OqIGjZGcWtKY
aRrskJQbNuA4xxVXv9ECjC8stosXUQNFs9ie7leGq17bLm0mdFGzLOI9K1GsUIqt6l+dO+iDSFH9
qSmKFVX9SILYAEPDue66LPCtY8wJ8nrh7vGzS4KQJcI/1KyCq+2nVf+4snbg/cc4j9OwXMXIJrWn
8XlA+oDH+6JcXJC4IXPBV2eWLZwSHfN/32utggdg8iL5NWAkiXAl78/o3p7VMy+L+Sf6BitW0YZ+
rTmS3Tn2XEs8vbpE2pmj/lwJYthaOWPVPR38Wmh8LGw2uPyEdV587flpzK/do0LmlvO1OaR+e8U7
xs/VeyiETmYHDzdsgMm/FgAoGuXo/F47sPJWUYLfaMshL9TX6Gu7tBEn/HFIs2qXXq0DxWyxrSjR
0LblZWCNN7nERnD6zVuTPDsF7S0R2AKWjNKfCRGQx5Ls9IBsKJlWfTwCHOIreDHnM6O2kSeucib7
IEy2xu8jxyP19LoohLjcooBZqslv2UyhwZXKfHNhieqKAgFCHStlvWjq6EgORe1ZS2Dsq5IaQiNM
yXY24QIYbsqXkEobuOQg02QAUIdBwzz0qUQx4D5+QFGR9qmi5yBScwq8AkzAedZJXNP9LU9cdXWP
OyZHlO0h0P/qeNKob2DggCRZoyp22Xa3fi4L4iHCNhl2rNSr00Vq0dZlxZZRLKBLQbAa+6d6fy7g
W8EKrdmesJxEwwG66PWcxhpyA/5KbYzDBFrIH1AEr7YEnsk08cNORUc9ffBOujH6JRV8yiroGMS2
iPxGnxjzhKR+hWISd2k9/QDry49xltE8l4bBzMUF7GWmdp1i3+eemmTBHmemcQTUubKG3JSvGFCC
4MTK/BFDwAx2JtQjix3xWaYMSkaQfJ+zV256Ihz95OoPqvw2Tvuo906J2J0ZFAQRaHToamuH89sq
9DyaiSnCZI4M53y+E6sfkbLkQ4Hnu+A67VYomCEW1psqTgxVqVnRkgTTReH+iiAydzAz62Mm2291
06ZBcrOoNFpLXuortOcGWBa2OzMesBPIPU7yNgewGaAOGKD717VDwUJbGLUdFv/jzjqMFh9cW+nN
kX4/vlDGV8+Mkr57B9F31PUciaPA5FSU7i7yIsJbCy/Uye8RkwwS3B78BXNiwdT7x30X23e4PP1p
Qk5YDsbwfGvkoOCYV3+oJixcz7WjT27wIcDXQ6Fv0Na5B5hKUmscdxMS4b1eV4RazHVNEraLM6SI
SMyJCVBWZdNI1BTX7jk6dctLmYyuJIWf657r1SUGnbbvl6tbyHRxiiQF2VUL11s4AHBVDDm2eRgT
bjZNyFoVLYaXFNA6GSFxxKh1ZDZa7OPNlMBAgiDHe5jCWCqk+B+toyL1gag5uvPnFOOdnQ8V/NMn
J0cev9tYuqwdEIhPGrL3tvJmwTOrdQouUN2xXw6PboLrQNev3SbfKjRO/fRivT1UrpvB1Nk0e7kh
tYEX5uzO3z073pLkX4BXQb9DHi00wGQ83qk0OcXmZrzjrsbevC0jULT9IowEakkUMoQ9XmQ1dVI5
q744pLvkavRdfJn4WqH3A5xyJ7ov8IUTSU0Lb7wDD3f0kMZc8IdRh1TCcUsChm3r843zif3Tfxv6
UvgJNyWyzmHtGswfE6LmzJyOJieKlXAVan38udAGTTGr1CDKhkBOZMrH5k8CMO2e+Tm1RQ9gPKo1
Q5ASxE/Plbu5u76XiJcJbXdgu/0vRKhYopO1RlqzwYx/7ksqDApBlTIpy1oZYpjRTqOABcRpsaoE
j8PXyizwkZ25XnNPQp8CDlGMPva/IEdSwU+cL+B0xBOanO9fwECshURC/eNl43xwpkQMnb2225zY
W2GzEnged1KwfZjRZSWDWZJQ1+/qLOmcd5t0bpMslzWiTygAohNGdE6wwWbqM2227ZgBPuk1vurD
Xg/TyrcHiNDgXoE2ANjDU4FnO+PHFmm4QJwb00NirMVkC/GXjBbNsLnw4CTvTs5oDU7cIy91H2CZ
qPXJIawvJojVLjLQFiumZGueW/jSoktmbGTj4j1wcxGRukM9VedwmTukDntx1wndpB/fyBsHP5MT
ksW3ow+FNopZvbwo1dXZfW2eNrPnk4VhrbMhJbITi5rWeV6CgD0RWjQzQF/aNc2wQzvikITrlvsc
+O4SSJrPdjy3vlCTLVkJHWog8DRc7QseVcEqxIqEX3vAa1F/I5OmCPwpRP9e2oxUrIZJo8Rz1Fhf
8qQjahOee07zVB7yVNMNTlROAD7Z3T/z9YkinAMKUW6tdC+bcl2jzK4jWwyEaSJRnOlRb8HRmDxg
8upZMbr9HL4+tUCoBJp7OZlEQ5ZwO0yqGd8j+a1Xa2rNG+6YI+yI7a0aHkWI9LH1XSZPeiOprf+d
sXh6vIGwMaxYlQzUJ4LO+XhJB2ItbHGOf2DIt3ir7904QD8FbtdU52Qu9KbTTJDcM2N1HGYk+p4j
5ePdZXdZmES67i+VKiasqMvcBdtn6CpSQyxnfqWaETzA0P8Wm7sBIxEMIvO+Dw+3vdADceAL9Qqj
xX/mOqmsjT6WaFDft4miO9yQ72Bv+M0W/eTjcqcpKg+LhGh86PcjxbOTmNPDBgclB9NUYV6gtNDX
nZJBOT4VbF7oOWuHklWzkhWbXr3OlkDY4zzgWIl4FukrS+k3mg4UUhDUkv+oLTo6Cu1LwREYjywr
fEzdHDRmzDdF08lk3mbH81QrMDR/VX1zrm+CniUM99RLrJXjk1xIT8QTAnLiUj+jF+/xmlTPTlHp
/p/lQLqYCQwcxEfp4h7rmEsVj4j5Od+aTlBD3NvKqP1RrlIGhXhaZxGfT1TwJyRjuPQ3hQGYjHaq
vBUBctFZFlbeVyEeAXB89ycj4Ta1nuq22+yUnTNbsXtEJEF+hFOCFcpRQRi7P4udvbslVJORTIjc
3vrf+jwfmJc+m4numqPrMRRsxnhqLyjb+YZX7YLUCuJXYj/uiBLzm0WDYTfsvWYsrr5NZS8J4ll+
rRmEmoOa5+Hat+pruGtV2dJhbeFeLpK9zD4V3f27ujv8+wGVwe1PbrnuaU2LWpHh5rDw+zoJpduO
GTudBtDhI0UrzK6u8RQtzn93JMoq/MjN1ATvDMm/81LMQC02kxl7S/veIIHXfIWSeN24zxYiBd3I
2uoU24R2GOgFwhnU0zmTg0ln8eERxCsZUhtrXEtADhHYt8vY9iTXvYkRqQ1BIN2lZvcALjwsZ4qd
OgsFJrEvGuzHqukUr6SoYCycx7DgNvt3BDvjxFc5zMjiZo1mfdHeCx+WwdA+woCW/p2ZoNT4HeaS
yipQzaLIF/UK0+fvjpHF27HE7AIHHvPTGQyaXV16lJre9ayVosB3vJYE6Bv4TuAhj1ePEpdro9Ry
u+wYIc41sQ1Pd1G5XnDmNM4jUc5f6WOCucqm1/h6TceIuBjjGF7WrIOQR5zXy+oe9FEREkFATd/n
++x6tRg4EXOo1lzZhELo/1Zamq9WhaN5A+QMhuL5FgmcSlYMi8GpgPy+C1gA5YDeh0RBcZTSB5Xt
ionVx+vZPXvfPTIFqDDtKceFOs1Ry7ps3pK5N1B7/LM3Fd+fNiZXiQCO4zxFrTm48Df1aFvuVVVQ
eeHIF8P3qa8+4UEIknyd2OkMrKX1Borkck3NtjDfE284ZF5P65ZCMhQjoLYcIYViA/X0F1RHwoTC
u8/0ZGp/5xDEliGZVIZ+70H92dDT3/jdHzB7yrRFsBJjGqEGy8u4065oJwxs/EPp6LzUdAx7m/vm
seknbnty9b7PSurvwvcbnGhasePrjw2J8WL/sbMQXqjoAUAf9i9K4KaZJj8VzUlze0eJxW7f3xH8
89l3nqKxYSsEiYEC0TYILyo7zNSLcDDMXl03j3j/pSRKOlZY8FcliaY3ahGIhuecR/mKjt08cKfg
1sjcu5tun4EVuB1gXQ2628opkh1B7J8IYrxpxVucCM3eaEEn3mTJQCtq9k57uF1f9UYBggNS8YiD
qMHaRGote70S2jUjAT0oQNN1AU6tXBdWBRWhMGFZ21Bc28FOky7WF6yM3Th/XUXbgIwB8iRLIQJa
bpZxU+LdlFpO428D9ck3C9iOw/mk2ZH1XT2IlvxuKxXxBRSyvVlLRYiE2qYBwX8GoWMDLSnvH5xA
BDRttVEqV4uE6IbxyTderJ25shdiDoTLdT6ii9LeN9WnLn/ZjMW2IFx47SHi9sJx7mvW5JYzcVgh
OLITC9/hHTe/uCWnIU9SNRwCaq9cAA7yHz8nnR8YBke7ESMXFVSZeW7DwHTRfsXVOhxT53qpN0v0
M9l4482wQ2iWZlYAi+obCO5g42KDUHdwj2ATmcYoBTxthyeQEBLqQGvzd6s7K6IdZtpoLgWvRBNI
x0MHKwkvzaGnIK67Z/Vd9qzaGqBY+1LiPRijwv61Gpy4Y0yzWw/VZAap3qTVNZp0hIDOYXSKdukw
CuXpspOZjOJ2q+mAJRhYmutst0uEP57IYXSmck/Bw2sWet+wb516STx5g42jkghmosFm2kemihBM
ewOkiyHV9a/NDHq0loVYl0AmF0OmoTWaORbTxQEig+TWgGYcD/hmgTzxmnUrNNGg5C8izNDwy9hG
FyTOktAONxiFRSwWFF1Ms6Mj/Hemie7mEIv8IWI26pqr8iW+30tbdl42ORPA4V5LrK3VtIRfuLIL
CtVFAirSlDj5Qq+5h5vbkOzK3d5MJsJwmLGVg/9o0NLsGn/e61Oav/hGMgFwGYynG2mMrzHOHVrz
3qCJfl0JepkPOmysbZJuZJ0uilEkCzZ3Cy+jJg3Mb3/lzIv9I5jgHbvhq16zQtt4BR66F3V6V2c6
vll5k0UpkbktWcO0MOkl7ohD0xdyWfrwr7mPjqjxBAEy7l8df2jnWuUdYKcUZN1+j5bsjMsW4gkT
vpG/KYM1zDCzJf/0Acf4PwfLOevzxQrsCqUy8kZdSPKEDfOpNBbIL+BcMI6goEU1KrRNlmmhS/SX
gPWt9t8aDPV3jgarTlWa5M9/xRz6UC7Xddg/itdDwEtls0ij+7LJOQSJ24Y7Gwo1hc+p+G+4GzoH
lhioKeh3mCwP7QkbhKM0tcga0aFI4QA5ZxxnnQ9iDPGU/QJK48e6QApQFbkCoG1Jto7aJUfDWtGE
Di1VjV52lD7M4TPCj2MmVv9HNbXOMgXDF1d08vwOnNXoVtxwMWIlcNTFW0W4DYh9Lkm/+tMc4j0u
PDhNK35wTHSQlis8BbX+U1Ayj8awBNfcdws6Un89HuEFvEo6Rzvq6ivVx/aoHI2fTVT9qa+BiNUS
5VY0g/B4u0m9tNSAbPXdW1yTncYqh4SH2Fn9MjwgvV3otJcWoVKdZdyERWz33MJHDZcZYD1rboyE
SjvYwDU0/90GS5sAytL314BrsXB+QPt/IyFdDb1BlT/L4E2KJmLyHIMPFkKCm/f8OjVNBB/2BCAM
cu+cWHS4H/8YUgmWG1G0HY8Y7z7A9OpqdZ5/i5RK42ezzxhcrFYL0H+0xfvYAInQa2wVGgRvM37T
8NnkuQKIQKYYBakjOBrE4n5cXAfejoVpPb1KZ7OZW4gK2r+q1GiaUQuy3c+f5d58ztnaxtQuTX/k
aNFZh8hDWuuzUcmcOajWRzMi1yn++dRrfkgmNLpvON1Rbrh91E3PShg4Vyvls5V1UyVzvG0jmGM5
TnWcbZMFLn3l+iZgnZYDsvflEUldbpaiB8BOXpjKUPyWapQFfdOIP9SPILj0KIt+/u3pIg3C15oS
1xExZioZirbOTOP/BRtI3hHRa99Omn0CmdYskUZtMv1fNyerPXL+Jm+ueT3yGElsaEpxb5G9bUtK
I6WaUBrTcHFy6mg4TloEOA1qFgn+duUJ/tJBE6CPVWugIZ9YoinYjF6C4yEPzbcYbhxgzmYfmWxu
PTugKNGIiQSADl0zX7SEt32h2C7+kep9hKZ/maUK/6WBqTRUuPoVypfnjjkO87e5cdXCfVszNp41
Yq9e3Vqlr1R3aDUnT+tU1NGF6PLxKWBlE2igHCTpXGPc6W25hGy4QQr2ST2MpqrwVLKH8rAWmW8h
bVCDEw9wJlRBuo+p959ITAtTfCOSkwX3WzIGdMRj6hg5SLYDpogQeEBnQ0N3mZBb/lNQhXMDDlll
4zYdVJDgwzAkuSUSxuf6mn1ev0Pvcep6doxm2F2ZejtwrauYW9DIANUhvPfhSQvbmpkqBCSYN0Ao
MeAIJYE/hgFzhfm1AIbEacAPg2omgOQNzlNfpA/0hY58uDRkx1XLdZMGhn47grHAFy64lbhcv0hY
u6miKqUTMmtEH3MCi2BjGJOBroWkFatfLpH4VIJBvDojVpn97eH8XoxuZ3oivgOe8jpMY4WLdb/S
wLVEEGS/1hI8N3xdSF63S3hY3Ndz6POQeVfvMTZxwNsyPR38/bUfp2szFqiT6odlYwfrDNvAdIFX
xT9e0IiZgdDZsCHS5fkJZhB6sa1welhDtlPP4Sj1uRJNSslBCVaIloJatHawRr/iiRZqZhk7N0xp
w5uYP7XVzDmnv5jT19kqM9Yx0fsgzpEeTjBMj1Y1KgS898I0k+3vdRbiM5Kf48kCg8eXW6Zaa4Uf
v+VmzLAMc6deRDq29mezsFq0a3zGwQLI2+3PIU67H0n1MCON6fSvQ3f385ORXX6v0RqmgqyN032N
DpCwZnL8yvxRC21K/re9OBtIFixLAk7BPWjOTH5t1LU7FgEWTWW4RZ+5s98yCvi9Jm1BuRZKEJlY
HTnBVa1qaxzpSQBlfpHfLqM4oPQGwClexniv81172NG4Ctw6vJabycFFc/nQpGsSrGQLf59LZHb1
eeQR5uuTHnaCpCo/yvm6sxYLvlAVP5LpGOZMPLuMt7Ew+0h/sywYRB7wQHSmHODgKfose7aX1Y1M
s00kv3LUMQnGFlOiV71pWChbJYKAcR/P3GF80GmgyPGOs3LqtWZygr8ty200kH2v4zmuxRsuRshB
ilX95hkpdmOPoX6mnomjkpKNL7rhAgEWP0JvIWUngFgSs7FCYYj7I77+ofh6WwboW4WrkCmuZxkg
rwpJMHDhkNks9X19nk13W1fQfFF8EiKim3TbgLBWrEMZSnHupg0VJKk5KtvWRfoxknnOKjL4jG+w
0JvJlOQwypEFm+HaDMrkcFDz8RBuy1WnRC3nIDtBqOliP53GoiMGBo5gCOdsIygwCZxm5T8V3XqD
ewS73Xz7J7UizXu0/VOdrLnT4z3e5s0vgGq1nAkQcBzDDP/Xw8fIrsykWn6YODJgxFhV0xcfa5M4
FfqdXd27xx1PO/TUtr8VBjhhSDrYbMyi0FAWbnGAKdpDFNyNpuz9W2XLNPf5rgtvgtpZmtjccvH0
lwUmmbn+YMLA9cLj31ElkbQj6ZW3Sv/qRoQl+1+9vJsCu+EbUrH1zVpFHrVc5FtyYaXyu6eXHBRe
mWb59lOEYkrT8YiGwWcn/6jx1O0oh8Am2yNkLYIILZIew3ZwmKW8K7bgiyPzMHaQ9KV8wxEOF7Uk
BjQkElexp37LYgvhTbym0l5ewTj6laNIqRvGs9ph9Y7W2ZQIK8yzMvmCVDdCJDTnOJyBoVHg6JxH
D7nP1TGe9x+fdu9pnTV/mtv/AnAdMRdmlL5fkNxlCNP/mWPzN4TP1MsnMAhlFaHE8WJjlr+H1+W0
iHsYcKdSzgH6orMeUu8J27TpN5KkeTICEA9E/WTbl/EGAO3PK+oaRnvgjPK3XUWCgJJHlF/3BRYf
EcPa856sJRCNsqGJYRslRvYLZQ8U3jgfnSpS8rDxOvBh8r7W8KK295kfhjb8jh1X91B33eHJyuFg
ZmKD3e9MBdtgrXnDKZLV9cGmbW7xjyRxu2OCtJakQFrq/K7YXrMlHZ0Jq0mqvNst1T25edX6Vuro
cNgig9FGC3BXMCjeKvggjj1wdZ1StwxchB1JbPQNk5D2wYGmf+8z4TNdnNsoloJd//JJejuyJM3w
L/qWwalPsXZ6g1M/DijLAMd4qJIMEqhEe6o/fT6Cyrf89TBjMmfWMB7xqDBdKqpLF7t4chVT7Knf
M+3HNqMQ4qKYAI0JnXm3Zxp5sFstcLMpk9n0cSYc9tOY00N0SU5Ew4WqtjsuDZZwIi+4XqD/xosJ
NLaRKpE5JL7KtVnurUkR9LDwqzVdB6p+VJ1DYXC17LKjo607swc2kaXlCwaTz/xnuza/tUATnoCZ
UW9T8x4x8kJMF66VBOGgQKmfwrqwxDHttg4ur0ljYNwPdVzgdSwgSEAdvWQ7AtmRGUBopXt1ulwi
YS+h2wyYsG9by7Tv5B4nhOo+jHeGWUhQZZug5R2c5WdCCx1Alp3vtComXwsdUhh6hM608RhfceQC
k6dN/PDRUu8tBRt9s/UYX2PT5doHETyQGJTUzUOHfVriJFsf9giOIKttecaShUkFX4YflhCQ8qaJ
xLPVffdzB2i3zTCrvdlVfqMwV7Af6pEB2MIj2BBQdCcbteckpsR3+qbrFiErMo/YCYBmK5fptcVo
P88TnwOJFsTaoAb5dbEMA8kcJQtdNoJoCnqZiw8g5iSvXjq1d+nkf2eYVUdxWNj7FDfZIgz6VTDQ
dJy9BuX60Iv6Cl/Q5xdfTWNd31GThbuFuh4MCeck/ETmylOuEf1HEO7erO9cNK5mOal6kv4ufsPb
H9v1cf0r9xJaVYd+O2ZMTFWYSpc7dxi0SgJYTe/0GYs8+CqaIvKWDxTanpudp7sf4KqA98un/1+g
GtOtywr3rvr3E3X2Q80W3u/JtdPwBxjOLkPPDQIgTFP+CdXyhCWst/7Ilw46x1Uo/U8tjnl7Pe8D
HqhxkbZuS5FfM7ZleBlqjDPRHYIIF08szh9jninuWMnk3hkc7NHVLvfFv2cb4KeF8yIf+IQTmCWi
VxFcE/iwrfvfqr9gS4E6Xw2Gvr7M7udkWx9RBKyQq9GQRe8INEmEgpKmtWTUzvghiEmic6xNrCm7
KfVxRKAClrW0Yh7GDGpvsg3nI1rkPJT0rzGirmRS8uHIjvMFyRS9jIBRlI8D2f/Sp8BLlk9kWKtb
IrPgCcOiwLSTIKKrx8/9siDG6qbwXOTubjoiAR2/o8xubg123G89apiB6qTIX7uRGQxc72VyNBCz
vweT06njrvk8n/Z9s0/B+t15Vo2qt9h71edFHmYHQtshwRK/3GPVWkLar8ezGW+Za5xN1udaZoVT
k5cUdRAQNgOmlOJ69PtGFQRsxLh7tDb2xYgVrINMrimMtLUiSS/28wKE2UGnmw86xvlg7GLEhdBh
gZAiDCQj4EiMW+DZBzjJr5GKeWh1uLA1tduZbqR7XkFeVEBrcRWqiHKvhTDmktG72Fmsr9xI7FhT
PcKSDOQA3H7XMp4JKQXl6q+918i7SmIseWXeKLhJGERMKOXjNTRa9/pUtajMHUPHKlD/6FtoEk3a
y2/jCvn2xXRXuxSMlTQdEcBhRUxI8giPp/Kpc4DqB8cjVjf6dfLHISGrfErtTv0xA39uevifLt5i
mNbZtNx3z4mNEjSbGxLPVPycRuoZjtMPWYAkxh62deSKcbyJqjIpQB4XP15x7rBNihqVE17PPHXo
XYiQIPwV3VZsgkQxvhZLy2KsNmzzBoiuQB9R8qNjGrC46HqjEjVPM13+h5lBh9UqEXVVPoe0TF1b
iX88hoMaAypoc+jhIa54BTC4HTVO0Ce3wZk7gYW3p0fWxxZpgIOovU0BMSh+HQVdEj3aIl8++IUK
3mc9JO92iG9yGJbCiFxjnW1CojxfTAQarKIB7GH+1QB8ZvkWPK+kTcDlv03cnMo/5AXJ+DK/RJxg
kdP5jrQYWahWZ60029sB4n2xzvlq/qcP/+Z93vdJdqVvM01m8E1BL/v7hrFlgt4CCXDXYKf5Ns4y
tr++b9HUXfTpNyuha9i8s27Rt5r6ppBewsqqkp4hx3yEOk+Vn6nbN39XlIDFaYMdNzi/oNSdauGP
MIGomOJgmyu65UK4eResv85RqomsETWzLkG0OrnC6j/PYOFivyoIPYc/oblduNAA6pZXKTe15hSq
VlDu5OKUpFXnbOVj2UKVGuAyaGX46KieXy9le+dBHOzelNSobZsx8bh8CtkwHAF1bhdV8Bv0Ozco
vrC1ne/FBcQ1jQVMOgqKnXIZq7FDeub0W4psjKar8EvhF5dyjBtfhayjZupUMj7IG53SZn6LjaGf
b+prJQvtEL7W+71sfe3wkI0HejHgtOFqabXukk+FoONqF2kzdW3LpkHEnG3qCfzG0zaxfYHmoWpC
eV51wdiwOeNGLUMgbo+AEfN4gvhYSOd9wZKTaN4D/tLtZCAfUHm2lunMBiyHcMpnB9r96pmeMKrs
CtJ7Yj/XSmh+gDEL13LDYTKUpr12bv1dKcAPFUszMFCDG0+rgci/NUfgWR97rl8gt+obXm3plHoD
kNDpvS6+WXTxm/JMxlA8B4C7H0F7Uss5BHTktfeD1psFvHx/6Ir/GerLEOyw9YSJ8wtdL3ruSMPj
CncIC1gWnSou1U2A/Tn8GlanG5Z9NPgAchlaE+eXxEufjTswAzJFjuTFsEDlulOg1wpZ70v4BSfp
RrtwPT74pmTYmo31D/sHvkJZgfJ/KsOzUMKL+Pd7hiCKrsROYPReue43SeSLyyZU4DRlc01u/5KK
ntgfhQuEUd13/BkoLfz1z26fbdVXw5lvX1tkgU87Xyx7IESzqvZQWSj4WiWO48BgFVbx0QiA+mJ4
NmfOcmCfBVQq7KkXptNueMh33IrMJUkMvuq+HLDx7uaQw8wRrIuAA9ESjhEXfmSHNtsDe9/rT1Mw
AgD4QatZvBG4j+J7DGt7e9ou/B68qQqpa4AYeh/c8FDZpEvC38U1jVwVhxtDauUJzk31tND1k8Y+
pBv2ZYDit2NaQ9INvbD3hY8MFKsO+j4gN43HZqAMBc6ZnRqvEwu3EEvtn7Kmc5F4KV+L0zhMhKK9
zCuLF6WW6PiVD4l3O56dS5vZWg1i6ZeWnaFcVX6N3jeWfo10gx7ldUUmiJCxszZouHQdflSWrCRT
AQX8/OYn3bCFd5XqfFghVj332YwYIHgkhIzMGaGcIMCR3haaJx4fPqV7HnYBs/MrQzQjfNUIsNMU
M4rfUwGzlNLUoN2udK+513NPPEIQArs+6ektFaSPpn5IewndiSZinOFv0wBZFghfLkdux+JKCiQC
OMhVXtKYNSA8n32QFhqfB782G0uVbXzNKPcVUCiGFTdmJsv/HT7NnAFpF/LDhph9VFEaGnvZ2iwS
zOD7UQERZuDz/kMll7/JLDhoQFQm6Df9t9NpybTr+TXmLw6yIYNVROtkxWELzY5RYmkSJBvd1GP5
1eyrs9nnzpcmm3T/vKx7txDdYjFAlvvJ60Bq15jS0j86oLbYtWKDD7dhgEsexORhYjDNavkzIjI4
3GIqLWCWz0Tw9fZ0dHDkVQPBmuIx6QbmfYl8DJA7cLDM2XZR0rEmy1qIISqODS4D3s/VoH1ii0+M
fLu39qdpAcgeE3ax8PKRhj18Yp3qsV85rXRBkcmYUmrwQzz8ZqTeQIL8QhDxe2wE7j6KlBVJHULR
k6ky222zPd7W2b61K74j0TJZBW/ZkgbNrjip2nKYn6+cN2jqwSTjrev/25W9pkR97U4YHHcGU9Sd
WMMKa2my3NlFMBbbqBesEhUh46Qdv1xDRp0lV3imgvDyOPcj7o+QVIP9X7C+k9EJZpLg9ZeMbIa8
7ag73Vu0IDAj3XjifqrBm3bOecOv7r2eJqMptyGDB2wCUeK0whXI7HGoYZsc+1JUePvJ991E5zuc
tMvUq9cHluzsfjyd1pFsQwrOfoN9DWifJBYdY9Fw0kYR4wCfDQggjc5poJSlQIV4NJFtQ2vbrF7z
kKERq34TAs9bFMa4rnI60ARli0/MZQ9EmDwS/3Yr4kXtXZUm+z2qI0w82WbwNknU0c0tmrc1NYMK
3QpEb8PoJQfTFChUivMqIm0eEKwG4yRhBI++tkP8Uv7BX/BXRBG9+OihGjrwoH3MLPQPmM808lh8
ShviCQ0qBszIZtijWDJAYGlu2qEQ8fMLYyo0u6kEAy6LDb5ZrdDN/CzTSuYrno8XFJmTtqaQKV7W
btbfCAPuJGRIUYyohnIBPrvepOVmA5dj6bVb03WLJuUZB/q5P01Z8W/er0AyeOcv+59cnQ86bHP1
/8Pwf6Y1FBMeKziWckRZddKjYyX9vx2YwMnjoXLt4gBGDzpQy33HT14gPhIXD7zRYGuWiq8kcsw8
xwL9OFAp/TX7W9Y+FWhqtwFcrcKXQ0T7nLzeN7A3TZvI4ADlqY84SbFyglfjKGXRgparHPdxQa/v
PWxApkop0ufQje4537/1hqvP6ycBPcFvrnTM+Gy5UBX36eUv8RqNXk+ytb4xgZ5WyDXwOL7+6/bt
HkVYckWj/PB0JpH72HqQb7j08JDehY8wGpMO5xds4rptigiTyaqdI30p4x4DueqdMnC84C0USBQy
9gLNZTxzFIXVK8z6iuEApy/k95R73Mzs2VjOywsH75OlhukDjKnoLRLEtRiBX8qELozvJ+euqXZV
FJt9RBpJpGdGRvSI/hJN/TrOlN93L9dhW5M+CF1rmqO2VDrYfk8OLi7FjN/DU5QRFEfmcfp1EKIk
Igfe7iYQ3M7HMO+Q3HB38tjWD0pW1qMp2IF4NIyEhZisrbEkCw0z0W1j73PWy/xSIE31GiwvaDps
Xn9HfCQQ6tzrBE1ra9/2k/fWhYT8GV0nOX5D3ApTNewG24xJCsyEHHeiX6YGKxqVWOmiKBLYtTXP
rkVvChvLbVw+d1D/hd2MNyfXEOXjdgOm/ADLFtuC5ZBd1cWvu/T/rZbGWdH94nmUgBQXZe1ZXiXe
J5bWyhriYO9q56yfERH3hg2mbdTQzuuE/hl5WnHYbFmIdgFZGn53+w0jMo4x6GLITAKNjwcmjon5
V71e1Uc/KkGetG5IHfLfIh5abi36vWmJVkItxGdWMGws0Y9ahU3Pk4dtCfJGBSllruGP4x3Wknn0
prbivoD61C1M003LUDR+54PkYj097gm82DyAYDV+5+HqbiPLVeXDbduIzRd37jSx4Leoyqx764xq
51pnnQrvU35CoYr0q1M7Syood/2I3I8oP/9XZsMjSh1YRJmPehhmMY5nsL+SYipMecBHYfU9D4fm
j1f87anRBEuIyUBA5pFctkrSa6poLWxB7vDVA6SwhPxds39mLTXrosTV8jZfqZCUMNHqcwr87Bqz
ViDHEr7oAqaby6w7bIERMclwj/s045929nTtAiyKK4r6xNW9T2zSgU2rYnglouxAfLG8n9HqnXV7
wGMebaSOGdBGpjY8D16JZg7NMPSWsCPKV+47/O+V2fIIXqJYcZC1B1NQ90M6vDC3GQz/7W80K0AB
Mz4uPfqih969X8yt1v8lJHOcgteDqeMf5JAdc1hQjdpqNs8Sx4wtMrAI/0Roxl8SWO6j1XyuBGgK
R+I0jJuM2zU5rpoxCtJYd6HmyvVNwcKBA/upBQJ+ZHfDGHL3McKaMBTRV7I53rRPQkNJPATWP2dW
Xi4HvtoMKseFOawLLYs/xI5KE+ll9jiN/JwKg5eqO+tTcZaNskV8SHA8RzGLOYvxaQ98XgIUPMa7
zIReimxgY8C6PmCbyRJ3lOtCVuY3GJoSab6Auf/ZlHvEe4qTNRvst2+D7eoNwnlG/7T3AluJbCVd
rZ9fFD6LiK1dhmPatK8KIi23aMNUvkeuYUhyOgBiUJuXSgcp+NwvqF/+G38+urspQXARUYZaCZnN
qBXweIog8Wk73QLKeuCf/egcGkiKg7lCqDaqHVvE9eo6kLPAmMkKEIXdujZcgZYnjM3fRGivt4aW
PhqMRTcVByIyrjBsBSerni2azp8PIsomyKQyAXqEaJkPPfOVf2I7Sp+N9PUQuvHyesog6/Q1i9mM
1SpdZnyQ5qGGuJyGnabGdWgKBKBnX0fFKrMBLmcfnUt27mV++/rSaB5WVBKDv1g1pRYfA+mLolrD
sQPlTqbBt4fSxlYJqOpKMEb8AFldZL9RQWQaE0twz+qvV1UEbrFj4AQJRZcvTgW6PP9fqrpduGmp
jarn9krZpdE3aGJl5dO6Ud6L4rCwOHk4KGvzbIFrsYomg+sIbwfzVugAs94Wzxpaj2riuHUDusep
uI4NoGty6QeiQA/UtUYxC+S3wPNbjy11U08ax8FDBbOQ3Ef6gVDORIrtJTIS/7oG1yXRHr4ecK/b
+Zp8QkuOc2uSSq5dDdsTMFCQfugO+srXdjXqdUteGO9gjZMhisSTuQAJY1feJ65bKSsVl59IEd4q
KNqMRh38ZE4dA2ii1EXL1dYr3HOSgIzRRPVEw8I/WEWTXhVDZRNgXACGgJDSbfssOdBp5+XsYYNp
CtT0hD2AbdqptGYwZ4PTtIrkMllqfDRppIxwgZdBrwjG2oruwrTCD+W9Z/vQVayh1mSUXdUoRVFt
ON6LMaGGX3c4ze0Dnk3Z1BamlosreBOSEbrEQJtjGrebXF/dRre+zOZpu5zwP8fWCLBMZYyP9h/1
hRs3Ly553/tWMFTAh7nf9lu2GN43jFjk1PYIb6oMzsQ5RX3E6uUNTzH6g71cEm+cfomiIAIA0kdW
dakPanBpmNto3bZA6oTX6ozzh0cc0John8uRBA/HKBM10MOQC8a3HgIqZE8Al8yvDx6axV40o8Pm
N5VobqZPwabEBR9evT+treS9QIr1iplscIgu/aiqPy4GcPfHViWuUb3MFtovE4ObMQ1dmGR1Evrk
TzH+jAKVMCw6mWd5KPnMI9e910+wawaQjcO2t+vNkrJV9VJsc+G2MSi5TINGd99+yQA/Gyxf3269
EIuCwdr5rNkItzRh3xP1JYlvvieGDTP9k7UIuGyRykamzCAfwQ9eUuddTZ75GOD66Tdmnh/hfZ/4
ns8lywkXI0Ex01Kqion7yfbr2zwwk1JpA0ET20AduKBkfLau4pFMOfR4FF2BFsN9qeR8ccj402cZ
1I5Z/iOV4L4db+KZSg6XMA9lkNawqZImW2+rBsAkhnJvgVdief2TPSgcp7fvNaqilAwbXds8qb4T
ysgAvJYh4w2uorgm+B2CCiIhgHe7CJv7nIcqbeNBMfdVG2tNBKTs1Q+jljzjt01NzxRg1D6WX/YU
L6tCfo3IsE0tgJzuJMqatJFYi2EYEg2AE1I80q34iTiQ108S8tr0Vri3hL6MfFh8cVz3G0UyCQfo
yfiZ7qQjlbqtl46BcvYgSIz6dr7P0ZUc7xBvPysQxJ6WCf8mkYY/h3vRHkhp1+ZWIxSmQAnBrzCt
J2+4opCS9eyLJAUKmYk81JT0EgayGXho83S5b9A5QQ31IW6my8eEiMzCTAx3tKpbjWNmlTgObcYW
PI+2+0ybh41tVjf2zpg7kaQt05pSyH2AeDomTSC95iRCpyiv/Azei6MyGI82G/9dclKbjGCKOvle
5L8Aw8LaAyZqE2V8HrrVB5IIZsQILppgilKCUqRMQdbYEvgTzkV8YEFAvOCQ1EODuOVirwvj+DoS
S1CIO85c/NxDAYkOf/m3/oBKxYT51imjAOlkD1lAcIdBP8SfABLL0AkEQLeFL1SeO/J/7v6Mirnj
kf9GKMm2M+8fRD/HRVPkxmD0/0gWX4EF7fy7wp095AGBv0LF3iz6gpc6STvCp4CT3En7GI7KRcBb
SaWtFC16Jo5PjOqMJGg4EwoSjNL+lPpKzYJwkicQWax2D7VZZQSBfoEt1Xf/ArSn9X2hE01SJmMQ
pVGe6E+uy5UMbM4622eMwnVF6Ws19kIMVOf6yxK+ItdGFF7JYetcBlyMKGP9o+iBNcLZ6l/TYAVg
eyleYY87QUnKpuk+5pyVidPP8+iAKhKncURCQUmf6+Ab6lS7lMyF56kTNbTSO+x+78G8M+Vvp5Gv
3sLFIGVOqb4ug9oZzVkFocYY41CyZCTsAvGFsH4YGrBx+Gf6aOT+K2CTMmisDLuBaAzOUKtu2AVL
CclpM6pnotphRQq25oT6n0IuIhdnZBeHv8iIQMloBifJHgSW1bwBnqgcfPLJgBsBtxp5V2n0GcQM
ePIkQGAnvh6mHg39NAulmVHfdUgsDVOopCubpnqvVxdFYg7etBFu6Nnu4ASrgbulQH0TFWPvk0hG
WF2q65yYueRpschb9IeOd2J862Yii616UlakGVqE5AWHNI+aq75EgwND3xtpVtExQaD6nKy5wLcM
FIsoWfiTIQ4r+pR5E+HSMoY2iTxtRTjVfGwPlp7mMh35eU/bj7CjsxBDL2W30OEH2640w9AFD+he
5kAnk/flt3AcsG38XhSp1O6Mc2EQlHoi2N7budsejjGSAN43XdLMEKsJdoXJNFBbrQVulH8LN7Ff
goQ8SuJXzz3yE4VSji1LnOY0CAFDJVr0ZFVH4+bgTjJZLEvBgC2oBBGZPKYgTrnP0Ns4DutY7TBa
NB4r0BE5PMdkkKi3/GHPVa9Iut+2T3aV5uVOR9lBcxRbAu5+u1A5zf+WaF6+K/KVyD2vd20Bg1BQ
N6NsJ1kglgX422R95vMyHCGQPCRL5aA0W1oVEKbM0rTvNohnWul5UWwcSXhFRUW8p6v7shyUlq+0
cOa/VooeRARWyMb7M0Ow6ECNykdoTLGI2JP8fhoklS7AvuMMGRviXI+JGwZB0As8bgyqesv838wf
60sSEl7L2yu7hVH/ZThK+YXEhVSVgjMtW+q0r0kqZo78IOmP8MxokQ+MrbNmnijk+5OtQjI6Ngrp
38DUi3IVP7nIR78zTVKmiADP/aRlMRokes58x0wGixChs+bn9b+qx3RhqUsxE4GLgxGXpO8mnvjU
WEOMSYP0G5zWGSM/1N8Dzxcg8fY8yA0Yi4Hg8cP2XOtgcY3L7/T7GTaRP+FH95/H9XUpUHMQiMZu
/yMqHfYwIrVq+b4jqCcLKBruyERO+Nqqyg3YF+pT4fDi9qBNzitBaN2BGYch0hSdsuyul76Yrjyi
KLWjIxp8g/MzMkL3iG2z9AjE8YyhuvTghCYqWw2Uhfe6JdjaUcBo0TeSAS8GUhV57jkgHdIv7K9S
wdNfWrZD4fwTnuJh8xvNmoD1aaG4CKIimn8sMKKlsW24d7JyBuQG+8wIbdTmrWVlxiwFy3n3TVHe
mnu4xTEXdCNw+skCkhmj0WkTWWsIT8L/3TiwQof7/C2PbwChcnD2M2u0gBPHxxzfMmvqCT40wI5h
kJJ0MSQqD1Kksw6SJcN5gk89hqOISkJToVZiqBPuP+hWinQT7gK0Oc46/eD6QsdfuXciCZQp6Fu1
kHC2gywcxaK/Q4HQCOb+7bffkesbAfMnJjgB4yEseeeeGThCxaTFbuDceTWrmd3WG+xJRCwsvMEq
RUo4iZq5ymG61fFQ4pkIxT5WWyyfUIU0zbWgVcKswJdyhugYohFisbW/V2IyaK7ruRJXOHE7k5+5
pmXssB0FKqLVElgCgxb9RdCEZaCFG9Xrul7bi/gVeVCfcZVkB1yAaUrKAdZfM7xmv9kE29CFAyfV
8EP3hz/bF5gz5i2u6mKCrE5TBcoHxpsR3pTVKZcye0Nhb45AYoZ/6/bLp4PunqcDbdXQ6USYm97e
3S4eQZes/PLCj8CbCpIh4zlU6pYtGj6UmW5KtwlGS95DR1AAzja2IJJ2UoOQeSvP6xL/Akb+xfTk
yjNVeLsmks7fTAgOliks/P/88ipx7iAce4zGR+JNZPJkEg8+7lunmfWSzIfWA3HuUuicwuNT9dMn
bQk3QuCsa7CLBmJxF1b4JA058HgDS/Z+rZV7+tdE6pZDymK3my5bleZ4hywWicjARYptIMhVh5UQ
Uwl0y1oFt1Bdp66zP7VZhd5KFkUSsIKb6FjlzoGCN95Dbgxcke7FRKPGgX3R54/e2DI7nYoCvv2L
21UAvc1GJQFpdXRNtUjyEFFVP7vfigm1+BTLgj8o3wd9TnSQo5mNZ9VLF9mC+9Y6zEPiBdM9AlYD
xwsD2Mk+PmethGSWJrQ2DBjSxjSR6k+FglsKfuJqOg7HEwAFIIBV2GMNJ4fh87Q5svLOqofxoB6z
AOFCCWEA28a2bYZuCwtP09CnUE3mdPUhUVmiRHQHsnDho6ygbd3VsEsayVuHhyKJuiJv+RTdJMy/
H7/M+aJezLqghqowdBDlWASJS20HIvHcNzhqxhfMfTUq8T7ff3QOR64A1LemHjpxWysNFTHXuHQB
X0AI/OiVEhyiGx3XEuCW/f96oYpW6VQaziMW9VjH+APx2W7e26W8HgdzcXNdhdEA5Okkncs8K1Jn
Ce2+KfVW1QQottqs5jx9YGgidYARx92LYnTu14CnHxIc5QTt8LPMVd/387R2z1IQHr72nRuCckSf
3JGpS/I9O7eJjGx/RE4v/1rec76yBOjx6/PnkLvksr7O4KcqyF3cLmUfo4qQy9jm8tOQ3xexpYVh
7qyUd5RKuHnoRPPzK/7P3RehlhWQIF9wSrnpZHJGPgbhkg1KgTA9rBBSmCM/uUpNdNFu1STFuwp1
Qne2Pl/z1wGpa3ovA6gUvZPfDE/mh5b9eN7RZ9pOKYmFx2Qd6y4kSvmEYR8atbjWojG1ULW49AM2
J1U4focSAmXF304jlfjZ/RkC1dH7PVq/GBPcjGpIOm1iQI6CsmuaKg0i+gUI+kxUi813ptL/hcU1
ysUb0YV7Zek/VKqf0hyQ2tZijS5cWIZOuDgPyG9c+o+D2Pjy5BFZ8xu4BOtwagHrviRamD6uLWXV
8Y6t0v4bju6LpMZiMPRFbXCSss+n9UCAzXw5CXd250GrPfrhAeV0qNeID5qmq46tK6ivVqHELFJb
IDBW2EuCkEebjAgMizGKraiBKUbXPkyIvT/Y9gkgh4VrPNt6wG0VC2wd5noQBMX/2sMt1L0qozVc
0fYVPS+M5yp1TjzuK1/lQlzAYpjuH1uO/msmH82cXZfzS0QaHrrn+pme8eBQ6ymqy3/dBGdp0sd7
oCtatN/iruAdLKAY/a9v6ONPkNu4wOhmyn3H+HBm0sPU2FG/iFJdy3XuZnKfeCu5cdGiFzsQQdeQ
npd5wuA80WQlN95Z7ncCniNglG4ubcBT1zTiG2ieyN/RUe31/n+BgU/+HoiSoeaSm98cpGeGAOiB
UVAaxbDyYrXJkKZNYuPDb8UPKhKHAEkvdNatuxNSVBjJ9a8m5xWvT66aQNvt1TH7ORbzJVOHgAoi
Jqho3n7xs5gWJtu6h0gcrnRFY8kohMQGuV7DLz/WWf0wBPlQxZucDIxHJ1LmX/Z3CBizlG2dBi70
XknAPhajbpfKgSFb/hNVJEPNfMBeamlTTXX69yoe2qZw6q9MlU2uflArnFP4cZHSfHyKLkX2vxDp
vc9mZj64ww2+Yy5jyItJvfkOWutQxvu13AAxCl+2j7s8axYcE9iBj0v2xtrRSG5YV+9VIJOZQVGU
O5zMbPkBtHGhgOac4FukQ9D4xlc4y1KAeRNJ2en8oxZ5edXRbh8FsFaxO5LYw8T5LMuwA1JVUkMT
2Go5U604lnOIKNw1uJtZqbI3UWkAk0TE58TOeO5ZkSodkQYvjWY+YF4fwPb/0Q5QOZmTM3kqEf4k
lNvSQpCyIF7xhybKmgGF0iyYeN8TZA5tpU67B325VyqauWmWfJSrHqsjHDC+cSE3BdmYy47UpBtc
C+2LosyOUlC7umbe/HKmYxAXiDKrkEnSKUjLE8GiArRM44tyRHfwdjGb5J4MwRljkcKEEYvgAsXv
BVPzOwZCFv8RB89n3dh/N2GYC1q60iA13LoVr0D0TCxV516eiK8JwSg0RcjmAdyN1X8tXwNy2irc
hIV77Tz1XvbAq/CazYSBSO0/EVsYQ1ucXWrxEO8akF+iY5EnAqgo478Mwmb4cV2kptf6XEwXypR4
boNl1Gv8Zgt2QBncNK0nYAgqXpAevEjS1gfNKl91+avsod6YCbpsZjfvKINt782tYEYjcWVIj0qW
7HLTpsQMnUB8R1eEttgLUa48kAZDoyOUrCM3De/hjn0LZ8neQK7/YuCrdGL5NVbVdLnXm2yBvr50
4GMp+a+Q0EIoAiuxs/tLFUhWPnCyUBhsLRBKwX7JK/qsYBhZctZkTRuqBMPwrBI9yHPDT+qiJU7U
C4HroJiDh49vlWhOXCArUOfuhQQ862FUbCSN1muYa8lbBqW7BpxgF5jos1KyBVUZTcwRTbYXNX0s
AZepDICex+PyKMrFt7q3dXEahCscGdBMzTgzamZgF0bMwX8lOtBeGQpuyVDy5KFQt9TY5DMuWk87
PFrExS+oKjj4COMqzOJV93IiHm3X11XKI6oEJAH5ilGKSAozGTeK7lEdadu/BXCUHG1Fjgzrv6iu
+yRccAp3c+8iSigkHln0p1I++woXpbMhVZO2GN2ijhiYCY2lPxZ+UmgeR0Kv7wc4AhDra9bPQIpb
C4zzRQl4JuXMXH+lGaXpGcm0fIW6On1QHEkHixBdkRsGMVrJkEZECm6lThnMqbaa9jlbPCK78Py4
9vGPrwEvvqVKGd+EIbluPKJsvWuYOsXrWqidas3x1v+x4z4BjevG8eFdKnVZoN5RzhP0Smh5M8an
/rrHNn3mBtiaIkj3W8gShXx7XmFv0Q2T58/I+ZsUH/J3o2aW53UkxJZq9Aee5BbkozgqERMns0jm
prhF3TrdSXi9rjCLWWYP69aFCQzhCNP0Tco3jOFUxTDkc4xxOvdkqJN6ikCLvje+yTBdWjinlDH5
gnR580weM2+Z2UAKerc63FEk4KRibWFsYrxHSe1vdP9JbVKjqYAvpJ0xL7z4E1MHUthsDpSCQPgD
wqscTZmFYj9+QKYwncjMR7hNkdO+DS5n0gLmqtkPgTkKSw4QAUdCu7UuF9yyKYVLgG1kOtNa52Cv
nmjj4cxoaextKQV5KXX15az+7Tz97a6bo0o5DBjTYYXaE+rv/dO8xalkYDpVL7jjzytzLwXapweW
AMZMTbEkiVyCk0ZM2EhdPL9S+2Z1ml+njuQPmUjbsZu7XqVPQUEyTSspCCy3Yl/VxSs6YLmqpCYw
ac4Lw+ZnlRWYSCk+92mX1IoEYLbxjWbCUT4UmMMdCw7AF0LUbJzngfrqUh20m1LPjiaLhgA6u1mM
MTPTQbym8+eWqT/n3sPzUkEuZ6YqYa7pfmDJtzKGLmPVXdH+tft/nKNd9Lvsw0glIwX9BqXBKtII
1N8xBMmtsDsDYWQEWQM4Ojl/a2FFP622ahF5XGX6GLimbTbbuZ8uJiNUB3ua1gTIPbQYvUmYEuSz
ZlIuO07u4my+hkQrvxHwWE4HL9nxu9QwabCQJVCjoVTfRg8Sk78JSjiLwkJ0805cEGF+9thDjnc7
nh7vKJyF6UP33ckcwV1hOQhQCMu950NKlN8CLhiLj9UDLMU3KEMIVm2rMBG9h27c7+yPFQ3FOyEB
UIkqbBxzZNrmLrGXp5UexjyTO8AqAqK85RDoJu890+yTPR/ce9sMf5Kyx/jGmJWtxwx+w7inGyw3
LZW4rTamQPZdufXjaOAN4HpqThbIzEzKU9RzOuzyCaBUHSmji7++9n9eVepkViBbc/UstVz6/nvn
bHMfU5344hKd+ix4aLpgfcCohiek/8HqCJ/f5so1NjW8f+XBrpvYEiGkNWQLAUQEjIDBxHMeanb8
iKE3qOMi62THXQrebDFsqxH0THpDQsHXwolO5jfQnFLW2/bmBdeNZvaTFy8VinXR4zG6Y+IZZXBp
ACKVVEUrDGB8RPoGdVUQPeY2jRLvFD+MVQAQ5XM3OeCa0Ehr3Q4b3iHWWcIrxJYIOY3g6ML3J5lk
VJGygCZqBz1yd3uWWA3pch5zvspWUqkZ5jsu7lGqT1AGeT7g0wwhx4WfD3JFdQlOueXfM4gFm7XF
auHLN3eLmEtlTTKwd5WKCI2qBp2bvvg6zCtC3TFOLPquNrqDEa11jyf5qhiYWv3e2/7BVrcjJJ90
X9LjddBkBtgfb+jL1CxOmMuKL5mf7UIoDBSXV+rCzHlaTEv95b3b1ka6umCOSl7qxOmr23eeWTEA
JbZ1PjcYnTrN2HT2JITkTDStWJUn3zFGhLD+s4N8arNK6heUt1bWbPnAGAzmSkTms6+412EbrLFV
GWuN4BJhjL1X0m1+xomCyh0skbueNZu1wwpvqSkUXL0L/Q1/6msPGWYsFTkaOq0rMZAoxSM1c+ZE
SiTFb3JZL7Gb4h5NrqP8xGfN0qTP0bOvxHIhZ8616chG+4evF6bQu3CtCxcMx94wT02IPXgKa8CD
has3b38fz3QspRn+Em3Q7FLXDCqeFaRD0X6rypoe2pOH2aDZpUbVEDmXE6gadDtXP9MEXz1xYnQs
zpfpyzBfwhQrpRF3bhe+5WRLdg7so0gE4k9oU2q33EXZ5mcMhfeFa8qL0LcCPdAld8xeDxt3C0yP
3JRCUm/CTs4U6xEvQjdXGvQmVonQ3K56fCBIPBZwWMuYe3u3Zz3wS8ZbIfUBBDadMMScvoz2o1Yz
cuZ+p1gODPUQUZhM3BbcSRdoXqAsz2tPFBH5L46UQrk2hzTDMF1uYy7Vczy7b64a5DdJDmX1zxRY
2QVWc0ZjEdVSKlaLA1/Av7JU1ye4CDhoD7oQq9UAu143EcRYb5jqn/UT7T3zkRZ+M9KEkWyIixF6
4pugwD+usuD9g9QEciZEEBXXC8WG/1ezw7J2sVKTPsN5m7hoEdS00DAFNrT1aaY8PCMsFSQwaBuK
d/w7xuUAyyCbaRoIhGG1uY7qu5RIvgT4RozMWbAIu3GpGqvDMuWe9cy13mw2lUT5qYDpWvxzHAQ4
tpwMT3W27GZ3K+ku3aYlYAJJgIRVR5WmMFaFALCP21INVPT2wiP4sRTc+jrziSNdVv8KU0is1IbR
KiuuAdzIOzeyEzx/DUTJo2kIcoJm0TATKRxG1r38cGDzTHuTK1YOdxtkdRHk25I6fNSLAipmt+X9
CIqALE8x/35Td2YgQKbL/nge1032+4k8hd05EwdYAyJAgi6VjTUjKt5bmEHJ8WXRbH8AEJeZuIMP
qBRDqs5wdB2sxhjNF3kZ2XN+zNHiHX2xneamfqxm6n/KEjJKLycGsvjydtd5kyUBgw9O1to02+EM
l1JopWMtvDjvGCyt6UQJMUOJyqF5TndTriq3wT/C9Mb57UBePwbUy2uSR8RL1YYbClkMyiCiSUHG
HP4zdMPgMvjCzmSLP7aYj1UXzNKzbn+6mDaJaaehrsY8tuo9Vibg2SJ6orBRvQrAZg0npZIoK4ae
LVAClX2wU7AxEQBhLsGgtiEHntxbxnaHYA48XG4iYAGVBdJ2BdgifHE/NXJ4aaxOdT6MaL5tWqss
qceU373qSn1FUzczf+CRptbhSN6Q4DFpwWtbJuj/AfkMjZY0B1m5beFfadRYTiG43HuE7lBamP9q
Y4kva41UHpCUoQ5Cm9xIN2DEuU4f/3wecNpuZ+xLymnC1M4swdzERLKI7zLTaltwgrZ7Oh9eH6Hc
wTIK70iCjjvqtRz8mTiKlgHG3FsX6dVgqmsK32z526XR8vBVK3xr9jQ9MwjbwTAczKOUhiEaCxhf
ItaFQoiImG2PdoXEnXxSQV2rKaOFuIbc/wSFqCgm1l7YwOLlXoLHJYGt4QU0JavIOfiz66mq2XpX
5yjPK6LW/0BdqsFOsxhe3AUwuov10zAgcnuNG7Eb5avttCMMXcfAj9QmZF10y+cbjAgCwgqLS7Vg
HAemDSSpUfj6fH5WusjL3ltNh071ariSnLJnDrdt9RjygpUGP5aWKERqnZ/w+xA4K7P5rPoY/ycQ
Wxs+Vd356Qk8L1pjgS+Y2SzUv2w1TqUclKHoj90eRuXbTVfmHcLWZH6/4tcPKbdlIDmw7SWH1P/K
wUI9YBx+6zlHBBgCryqBz1pcBO1Yo2x+onvrYa5I95nBRf2Y7wgtIa4D9c/1NgtT6fpTiWEcDdCB
uvZ0eJTC+ibwGqTXiWdtcJIrLJxh1w+IDI/qGRtoQnnHkeYF8d2mMcJ0WV1oOHL2Q3PhAZZTkT9X
25Q0oQo66chiJOWTPOXLiK17Dgoy7WIdiWykppxMHoFy3qg4S90r6SPorIohsDzW7TfxVh1GRhaY
zVKrVVBMlAQRFjRZt8f9xNastKtCrmqcPTAkkBwyGJB3bL+ZhYBN/AhHDY4rVqY54J2Yclq+xaII
gYNZNDTp7MpHHk6tq50Du7Z/Opv2mXOrz3QFv3GwdcZjjStk/wkWQ9g+LBx6un4vNURtYOtnZbOL
GLvrnPqOkoZRqGPXWnLXH7CZRGEdNUuYHaXwU2thet7pQaVQ/Vy1Rv/azPLUZFZFtA3ybdpo9H0Z
DPfV8v+3LcaTfcK5lMnzocBL9QwOS83AZEVMo4T/lf9jD/U9/VU+vk4RuO3fJer5IoM8Aq9A61em
EZAILzq28TxSEje/npuDL2pa3IQtZWqsvGDG6wlaOMRL8twSPwHktnUL8Us1cgRw2pT3fnYJp3rl
ICDt1sQcbXfUKVFxSq/Nev9s8CIMAul7IyEnZC57i9N5c9dMuAk0eDh/srF51Z5ifOtRb9IToq+v
+yRux08HPpyAmw1nIPUtrlFSorB67sGNM5GbgcvaDd3vB6HsN62vQ8tfn1wK4ittoGT/GRegYHVT
DfRC635vmfqY8RRWmJ/T1YTaWe5aYtQs4gwKiwcVXO7mzSjRXqXZnAt+4xGHosvAWE05fI9/+zmc
nbCkSy/HfKv80AFvDRY3MZlJ2XL6QzUwIV3O95BGcQFQkn3p0beHw7ZA3J4T8FoOR6tTw/3uTZUB
aaaUTU82AKEfqHbo0VoVnh2XWA1FS6X37D8KJnDEQzMXSQ3Rxu32YDZBX/VIR7hAC9HCHZ/MDVDe
bnA03qtI12zpPIxzIRMcU9G02hTbMMfRxa5D8x7ZPFJrfG0wT9OZy/f7WIE9SMeHKZiIA2Z5Lwce
+S0WXfpxfSMga+6v9ViUdc3RelEdNiI7Lt14K0kN3cAId7izQU5SL0jkf/+eJMBL9izHbDUgXTw3
JZHjEnOPISZYKSKtomj77buj6HbuN9CUUeP8ksmJerFfk3FpwRyFzTu2CewWe+vjlKiePqm16raY
MMRt3JhYlxQ8myILuhTSnYbfOBNX8LVcNAXeh+YuXNG2c2YT5wkj1noRc+EDaTCQBzwBT0d2kkAn
egEAkPISlYCoCWD7nzMyV28/+cDfc4xrK8D9rCUOLI1+yGO0h0tjZNimerCRgpanieFG3PsaVfWT
BqChzpMffrXdkxQ6zs2ep30IE6naJxqyE3OiVOI2zayKPRdX6/lu3cqd3v5dJapDJE8DDoRklLmv
ys4VrytWGVfwCBnEfHGeiRTK6yjROOW2Jiv+Cc1v0qKM8S98QdYtN9shUu524jUj7IDvvTB2W8Im
bam5wfusUURzG0osluRjdL6Q7Zle3P4Ztx5OGQECr+Lyg4dcsKbnzzj6FJVi+qfT3b0AbtA0mjkv
ypvNZHKVPnHu7i7M8E8veK0HJTpWHkmtdecNOURLJ13bxniT+viZ3veBRKh8ld2vEmU3r+vH5ZdI
1WsHLdPMQl995wsn+IejQyZKKAqVnP3+k5bPzCUZS6lyzLMz5UrTtB8IPOU2vZaEmhMaO0wn0zjj
AZIRqDP9n/7czqlv1gxNUiA3bdebAxPVFUG6iiOoa1ZvBxA3qYDiuYM1FTWW2+v39DUhsICOkBLn
CPShnA6PhZy+wYfAZ4R8gcAB6qQa/UjKJ0smbIfc42tF9UIqCTO2kmTLXEbK/Edy9Ic286vGN0CH
AXZ7oGQZE2VL8dvreDkG3dJav443dKJ2o4jilv8pnLPF+hIBSnNVxMW8UcTEtdKkxA44eAlyCjSY
JzRJ8Bo5ZK+BJFJtJyh3AGR246p1AIYBFtIZ1lzMDSWWE83xiqEhwRHFR7Y5qLf95VrCTnDAN6Xj
vebPIMytDRWLLihDigg+VEt7Yd6g9uEI1ns0dLsYWHsRZ9nckjyZjqHCsnARbaeez9eHLP0NuC15
FSmT/VVKRo5qJJgL+/J1xiUWJJzuZpDapaXRWxVOG68cOgVgncGMrgvjjFmT3/XVUI/MG/z/KpM5
BQH/awfaykmig8fvItdCN6dyGg87Zka3zWXT1mobTGg+d44l4efeKFdOzAjcfpNL5rwpDowVZW/i
TWX3Sf1EMNCl14DHT0j1YhdlxvtZPPHYQnhJKCBv8pmEcCOepftYGhSVRX1GB5nlvQIzHWv7dnTB
iy0htxZJ+5+9VhJ+SyQaXOwnpSaxC8nhoFU2avqAQKWAMgiVcw8bdHdi6aankZ851nZYPj52nR60
iu51kspVRdhgxmP24JsgBj7OcOXg+WQFrdv6za1U0xIn9CUbWydbyfh0uAKvHQcywWmSkBnXnnT3
1FXD1yTAxB5+7lFZ31vZwSvHyb5gURm6Ac9dYYdKxIyRw0NI1QaZ5TtptT7TKXjXJ7ORumijdogN
MPZ6/H3mWFwQ8TYK/PhaNU42E3mxxXFRvkO++6C7snXoTMbr14e3NNRQ6L9iaAD3tofkQV6ejgYv
uvI4g/APW9MPGOdrQG/FFEMaRPP7ZhqUR0OQyxgeeHGD+AVIu7ZPnssYYFHpFPdtedui2C9NMxHa
xFrp5+75cpEdszWyCYx1X/zHcbypwWuKlaYejliUzh3NmfbuYCgrIGBviwb7dTxSdwEHYIszmtLT
AYb5CVtjyQ85DKhVLfRdVlnZAZqPvg6elw00zM9ASh8ZaEIDkuTglJPoXqtbyYP2Scmdpjb3OY3W
/UWW54zWtoAaD3gpeJjh5BgpCeH+69ncpgQvBS7DP1bWwgO/Zt79nIZH1kVXWlurRACZfStmTGDs
Ko068I1qLUhf7wZCRLA5WHI/1FjKV5ctaDtIZfT5Pj3ozA7ugDihvBj3SftcCNdJkdzzxw/QvtoD
qCh7+LNW31wxy/Oxbpg7f/s6U9LYEe/M1ji6lcKcSWkoQD+e0fMpv2cCymeTvrHzLQkwvBVn3rR/
DMmFdHw/tT5u3icdwtgk6jLJcG8Cf6jF1UnFMfrHflnXwTd70E0753e4UbJN/6vJXu/1kD4RtHxy
V49mQFki58v8hhG4K7vAkfTkSGsdkYeTctGoSypOAMndOMrvmf6OS6f1xSJl+v7IlqZXusqi81js
GCuHZUXaZTNs83QC7nb5PY8JnBgR/1+Ojc5WoGZgerbqCkOioWcwkUltG40dcRqDDHnlgmJXrf+6
JRVJ+bt1dH6HI3OMcLlXtkJqFKSgZNXeQKsMhMah6L310eoifeHxQUnbm4k3eCfu4w7W8WglaHCH
8LuhLZq6FygXtcBhMr3RR65LzwDE4dQVe0WEEpn+KsZHLo+W86tlD3flT3aGXNmJclcsr4SuwHRo
rbZl+Gzm3fZqbVFDWUnOH+khSn8zx3YdwVjH+A+6Pz3W19KNKP/PUMLeC0PdPWOv9HgbxoM0ZxMM
IwUGvHF18F6zCidfF1dIIxWds/y6XfIR3oot9ruKizUVxV/BtppFjif+si+H3IHfW3UeOO7/VdPF
y407rz+0nA9PpL2dvlK+AyYcDDf1l7Ua5cm8YDKmkU8+O+bGLOhG/SIFa3pvdsu7VNjy+c40RpsR
p9x2mfV1HRThyHxzYABLCtKWMOgC8asLCkAm7Z4ncGfIvMd932RzK6GKqDCtzTU/HVVorZKD1Goo
wEKrjPpeHHblCjG2Y8vR12sidulQORMg7hmjIdbOHt2m0VMwtkCfmnfI0oexmFIM2HAPgvT2cXz+
wZ5FrlNpoaR1cpgWqkWyRRrFc5gA+5dZvfyCil5om4t97bV4Z0EERhtlxnbvm1Gs2ETeXbzphJDV
xmvkohtoCkXy/C14WqxtSpY6pBjk6lEPJCngjrWMCPDtCjDpREatj6sWHmy6EftAzBrW87dD/+m6
CUG/g0vO//gmqjaFasfs6GS114kIRdjqLnbYTFf7AlNMe7TESpREkjRefxGOUXTVezb9ESc/cc8I
e0yFbvwaAGsaCsr1i70qrUYehoyqJaoEObO59LX0U0J7r2q1+44UkQtwmogHf1UhN1KriWHBcYPG
mAyZFwrCIuDww9lidUMpklmdpypZBMJ8vIS+uFbfgN7OP6luqs+bUECbD3LfLMzOj9qXk3wuWVq3
tgtySZ60ELLu4g9WI9tU+soK9/shnRI0NQ300xa4S4zmDArC+ZGTAOM4y+CfFhGHiWa7QZTjIG4z
xOJMO4BvGoSvvAw/dSCWdgNmxvv136yfRGyRXX1lHSuVcHgF+FzVjEyPzdARxtKRbc0E1hWtOZYH
SVoDW8pCv7nRbzfAKf+WrYa6rGtAtWhaXeCBmvh8z/zmY5WIUQLH9UhHNUBtE8zboQymlaAHUxAC
aFSUvARHI1LXsNbHBLuszpABSpxxzBz6zFss77FDPy80r2B30JsREgvrJ5QsHHTGR+gIQwLy2uZ6
FabdvT3oueV0ZwGRH6nafUb0n72uDecR8NjwOjs7SDvC5QSg73tNjCAycGrWIyXgVLbiz35EoF5z
1e4jWo127wwwQgwgt0LRwfMNaXWiXVK+zIX+wqVTYX75OL5kb6xW8z8ZwWkLnHo7RJriEJ5l2oe6
F3hYUK9myWgT5JMJ7n7jKSQcxkDbY74TkItBLYLE0lJTNjQW4ggHUA0x84Grw8xNqn6e6YyO3wSj
IHtHi6vj6VMf2kC5z6SucXSAQf7LoGh+3fV/EMYMiharBx5pY0QoG7y6p96XjjzqHxh8K7g6Kk61
VCrhcCS9fmCL33Gd2a4lzc95HHVN0KubyL2kibP8u0z9opcre4b41oAF7LT3w7hjCB6Dve6xqAQK
OU5JNOBYkSLnbV+zKg4YAkP+fkhc7JwlXv1nMkL/ElpdSrXIo0pLd9LZtnWCJwE/+1gNog5DXZ01
H0Fb8+qzQrDZOyGC0FDEnqbp1LlDwDxd8+CtsugL7AA8aC5OOVSJIxB9autbjGfigPDqsg3k2np+
m0XAcBNVaz7h7D/oeT6vl0r9ZIoudR7XiEZKoxefNy6Hkq1E8oGr+2F1agfqSE+FOlnjQT+WtlRx
CDHy8FqJanX2tJ8Iw1qhYr2mqn7YifSd6QMTo01iDOrVPUgVmTF3/pCsAgZiGei8TniGhkoRLHBm
s7e6sAH83tOEWByGgPWgFF9IN1hlyhAkulUv5qPpiInq383hT6DzLaAftJMq3tG0aWIHNKMRCaro
DtOGpH5vsiuKy0A1hw75vLgwLZC7M9TsjFDJ+6NcKfmnAoUcffUiTm5+rTl5medSxU004XmzyuUH
R4Ky3Fu0cyKyY2dJHFPUp9KSji2sB/uYsrbpylke5FhnoZhpggESwQVxL6riLtMr8YrrVHDERAUg
q6y7LVcCKy1Y6oMdD0mF1DdHaG9rURoEfLXlk3GkcwWOtbbE4pPUOkwkiQjiVImzIsuSMUVmsdph
kgmZ8uxdYiXtqGmVzwPsyhPk5FW+o9YdDykOPjlmM3gFADSbpTzohwbybAH/jtLnNcnrTS2uZFDp
p88FUuyjUwxMKUKtOkCzRiz867kZ6ODdeQlvrAVhBcoaiMfkz0Lj+OjVDnF3zayB8jdjQJDGVF8E
jbyCdvRw0WY88JXQ7R7eEPCSgakH5IikH4/UChcg6LwSoQG1wpWS3ThILTsbS/xefYDtpmqAtVey
HPhDYXFATtOaVNrtDH2/OUMp173q3VUISh7rNDK8qu+0mew1yuGJpLvfR2WRxnl4EN65hWqCTd/M
rP1zU0CFYdMUrslwdK9JtEoAFd3RAnxQ2k5IZv6opQ0VBcRcp2Vb5mAHp/i/rw9r/fhemI6WCYGd
B/vYhJdrbFmZH/qDOXyyQWUNeAZO+6cZ6ZLzbjylLzzWEdNDP61WbgJeAVi6BFnl9qykNamajVtJ
awG2lmgHpegewof7txKk8qKcmlbLEyupbTQeYgrdiCwpoYzhIigrj/b8FyIYr1zGUF2iJx49zJ2o
gazxbHwtc6AN14I+RrSUmpF9H6RhxMM6ZcYSrU29y9jDKBuxIryoIXIVEfuWr+zk6QHd9Smopk5f
wABVB92h4dKIjkOj95R1gJYUcgFLPfE82e+xNs6e+SeSWXMd5kk143Ia/Y02Y3YtVco5XG5o33Qp
2N77GJkVrzwzlxh6ko5rMwSXPN+GUoVXYy3y5yBzUcakkahy69tm/NAQVEEcA6Ys5OYhct30aDh5
7oxgqUom7ZpnGWNY9lWfRMjBEgsKkOxkhyQtgqh4jo1JCMllQCrFSzXAu84g1hJBCZDWHNDPcZAo
Gp2khFVLpcUwSqiDpf0jSjVIjXJO/e8JvT/rQTtzT9SH2ACJYsMWjPHBpNfezQsb/1CXE4Y/C+Oj
VBzx5ylADbRVQf3o7LMbWSLEQYBQHifh0ghVAhok+bhlld15Cdwlps2LcwwkVsWXjQQMQOUNm1RP
O+XLT+PAeSqqig6rsMP15gbhk/gyEHyuFL3uOl6ojVsX4bIc1UzJaZJCSUqMyo4kAKTII8Siz63F
BKqpEoJzXKwjUvDBXDOE5ZC1LcAlk9/D+d4KZiLqjUFNjGcy1U71pKkQkINgHRpf1Z3onyTEcG1p
FU830+5r4hh9EsZZJtPpiptlj7MC+P6CQu/wy/HEoU9X7drskiiyMKKCj3q/Qc+JYiQEvTp27atZ
RRK5IQOnRBiapmXaSLbOthzc1o/J+O2TfqkU8ypSbuzlXbypaefMfB6BXVsvhyItqQA5mimt2LDb
PflctvDFHWbeKu/MRULqqb0kMaeuZ+JVPc+dpH+/OshmA/FidPzS4PzConmugYpdfngyEou1S+xV
U8Ifv1p9L3q+cYDGqJu7sovWdZFA11wzx7gIdkkMFVYsMpuZCBrdo6nJD1qm5hgPlZfG+XQN9IJ+
2gjc3qmqbYQW7boy3z6rwcdoxRrgnrQsjBHknXeIlSIxBTs3qgVdOAaXfFLp+En6zaeLKcBX3IY9
Rqe04RT8/2mbGazcaB8ZWES8ArkN841en9xqpxnfTwq2P3jWS3QHnN8xIEUr5/Yd4wl1YzHEP7Cf
QEBthCfvXWgwjFwzHflZiJJHj7CIfmznflu85QYU+D36HM92fjBjNJ1dPo0EaNTBnV1G57NouLk9
/uStYXdlp5G53piAwJJKEPnZpFezEzdLSlRVL/V76yHLOt/ldXZpMRR4StZA5+wQgplgd2PGpkPa
3eJWYV9fShqUTj13U0choizER0BNvJDTdRVyeWsLEfOnTZBxua0gLcj3EXNtSCy56sh4j3qlXc4t
y86umRwoz1JHKr+2AgIkqhmVDDU7U1+wzO5EVICwMDFN64HjNmTCbl5pgBiQFSesRcbk0MDoNzFP
UmjkuFfowjZ4i7sAxGgz6rDqP0P4rFdebhaannwENcBve3aVcebli7vNuga5tcubD8sPDKGp8RER
KMo3auxS/kF3EQiJkwFHx6fO3ZBLeSK7sz5e2jdIk2FmjaguDdGY7SFu92v+BbEgV9redW1ejnoU
OT/7aTEb7+/Z5Lzaq+4xrIxyCshEWCDFi4GJo76Y4xPIv1ze+Ep7GZi7CBJMGj5rInioE1Y85MsK
rmkomkeooY6Cx2HlhPeEvm2R2pmlS8j/mB4AJlCcwIxgybJUkSQmMC5X/fA9bhejy4bT3PNH7Et5
sVIaE9p+5NV9PUfQBXfU+x8867JUluoouqoq81gqvRW+dn+cDpeqG1gp/L93pMw8ul7Vk+qmonIz
M6E0qxKctNpH4/Id3BzmM+mu/F+PmkOAPv0oFFYTjV0l92aPjaRJe68zZVvWeXgENxF03ovhvBOW
YW/DCjnIGZeOKO+WtufABgZEaOtSmD+XmE71sdsfaeVdIxoPN8eYvMXyBjBdMZGGmkPSF3RICJ3M
O3tD69O7YUgV2prx7AiE4yRXPPm7HWEQL4PZvmAkmTWkyAEk4PopMgEEhwztBPXm6/JwyW7wbmuC
W/TZaRb1JLr/CLtTofnjY0965ettuZ0W4UUY02jzsCJQPGLEEBQmhxrG9ifQGpM2fzJKsPP9bC5l
TXkGsbP+JbDcwfMp4+9ISdB9x/wv6V5qQPda7LtkKCwZX2lXa+3YRGItZGn/CM7KTe0pHAZ4e/AI
T8y+myqc8jeHcPIJ2qTrfQZu5SSjiBiVbC+QGLiMl7MVjfIDkUn2WNnSwaAjZ5pHuIfLr/qYihtu
HxDbcYDXIdjIGrnolMk9kGydg1GmVUKzEvwIF5kxybt4MbVicaqQb+vU+ikGjM6XReUE9K+puX9d
8dsN9TIgXS1ydUwGff9y1g1r2lWjOl0Js5ufMQrjGtEsSzC0MMH10MTfNai0wPw4sP/Soyj5oe91
9J46abmDKhH76i766WFw2uxFjp1g3/fXGzPVk9VPiNyLpcgvd9yxRs2kXxwzs1YeK9IQx2BgftzS
Hic5zmxDAAQZBHNoSE45MQGnnt/AYFg2LjGc5zhTMyfwq1PtfbNL2/87qZup10XKI+t6ouWFliGS
a6qzB7s6MnOqT8EAe2puedFTNau5/i3HfjSkortUAm7HdtjB4HxSPXFrYqVKq45i4SOga5myhsMl
GRXHBYZTX2EGvgVtyiJB9F7wJ65/kVsr+oRQF90iPuQC0rAe4M1TArVCSTd5DMzaeHju02ZhNcd3
y7/FWH+VyBzvgaI1Hy/tKdXZJxSN8yzz9YdQn15wiZn9hoaTzDs3mrPorLVHJOqtLij7wcjsiQBK
XuSEDFHkEwCzuL/4NbdGZsx88c/kXLf/dKSJMLM+eBoBf/gCo4iK6uxCqj7jNhnF/s1o2UIlQNN9
ObjBu+c71/GdWPAnpfuZs8Ao82iVz2Toq5i0JXi9gBfxYx6uTc/xiivx9KZTtnWZCDxlUkX3coul
1MfB+BWWddDMAygK90VYCsz0u/cLhR4uZpbOIcBJeLUvINnaCd7Oo7Br9t2yxlK6IlAx39PR5fEH
5mXnFjvac91CJ61oc4AkcknIJotiI0oVDYrWGvjl6U/60OKOzlMlqcFvPbkxALz5/dr0PbjSiRrF
0VKRyZq/HcTbw8G8nv7FtX2LewuWjlydnzAPapl9SzqY8b9w9Xm+XeITko+W6ZUSCXpdQU5EIkdx
o1oyaTK9jXO2G2zA/ZzLBfhrMJN3iaw4i80KzePZxiFATzaTquHdVUJJ7G5BnUAphRVJDamylPZz
qyVvdz/uWMafjFuQDTyPfpIaZOJghvGn5opEtv9kZ0wqGqum22LqF4RlbdM2Ha1uSTF2BGr1HI1v
MAiSGvUgH0dtryOvUjZussGcpmxjEpdwh7u3BH0Hrvx+enbT9BsEvg1d2MsX92L+DfZWGQTdMPc6
/cxTFONqfAtNsomqOZA/cXBKInC2zFQ2BCkq91PDcANMu7il3xO1CdOejmQUwbTyqt4AzNcBa0iE
xWqHB1jaBgBop3iJsgFbTZI+KbxNaxGgUdSj3CWIWoqedYGtABwQphnK+dqJyLxaiNnoJR+AOui7
aeKD3Gn2NnixFgTGL0WkXGosoRLGwl+rJgsl6FVrYZnGjoLllTkRWvlgv03zsFgE0I472DWsDSGN
hnuyz10yCzG/n61G+QuQy/vkaJ6A7ddNF8tJ+/z3ikoxxpFW/vSN9/NCc5L/lCr06nCmEP1riNkh
vflzJzmxE0s+BG+4NAMPh2AW/PYa34Re1LFY8SDBz8Dok2q4HmMkCzCOzQcgKVlFX8NItJu45wGb
elhmV/CjuP2fR50lDq4IF4bHxx2J/r+qKghkWFvgfhDy8gqCdL+IQyE/aNEP3L/+ssG+yTO2TBQa
uQffFdu8i9tHoZQEN7JRbSov/vyzFpK9GB4yYwQqUf8lB3ZADVoUu0ry7l+YQV0om3T+VEIQJF1s
JJjKfL1WDYkzvBNAPo0tYi8PtQVRVnUHRDBOHyP7nLfdCE+sBMQcIUTajsOCjRXLw51HH8JvyaQ0
plzXChVmhuu5TVX/kWp4I89Schrg0c5nQLOa9PE5EOFCJWZOY4czYhiGNjo/ZVqTCPhdC8SmLsm4
uEVgRpyzjkCGwQ5tfl/Mzn9PcV9ismqoEW/44FFShOi7SwBFxOS6jorGUkkbYNoqquIQO02Keh4h
n8eG+Y5oQvQSgYY0rb7lBa+eV+x5PGMAw6m2eS7oKjlxEqzviETWm/FFjH4G32HaH7Z45fieHB6Q
25fcNbzAeUD1ukGO5ljstRLr6uJF3IOq/ptBJI2RatZVYs6YU7a6IUdSDwFFTFErLE/D7b0+y4e4
9t0lv/OrJws5pQ5/U7IJgG26kdJrC75zgEM/lx9sjlepIKNxigeHD3dUkbJk5jWdjDu+qNKCH4wY
8LbmCUZRZbfjh8HpCqd/kujv2Th6BPcByyui6Ez50GH+V39yrba5d/j7+kowbhO86MqTqMhnSw/Y
dN1MUp8PgN0Gl3mBbnTNNiid7u0fGKPoq98qNn3LxUBLDXF28YuMHQOR3ZOApP4MaoC7fQ30aI+5
mm1VACtSZihQ1e2TlOxarqM0XtcAM+j9fvIRZ/M68Rx6fJflCSVBWPqUfuxGu108oJXKV69RAQns
xJ2W+Dly917LCh8rGNMULDm9CJSqR55tkTOVREPnnhHY2If2iM0CfGqQlG8ziKu3DUuCaZCG/aOt
lwvux2WJkEzqK9z1Z75RGeXVMXQjukJnKlGBv3GYrfTWLdDg1bevSVEu59BFlGsFJqBzwJYdgrN0
BBOSMnOqM4KPoyPHGP6IU2q8liir5p9ma8dwdY+MTdJnZkyVpSOxLXONmBfp5ll+njNQYNc1FRIc
61PdQ0zQHea3PD9wIZvSEN/aANpgJR+WmSJJq3nXaVGX2PZvTY9HMR7FxSZv1mAKV4t/yb4/ysQ7
3wgQbp9LsIlMSOnKWs9sbEsYQnAoJaZz32tm1rfvx2s1o82BWZSFvIGX5NGbuKbMjlIdc2ARFPt9
M3GFImfeHHlInWsampIrClsTCoT38B5Wr5nOng2C6B9ufdUCQ8aiaxABZF5j8Y02MDyEQCw4NcmA
41Xv3ic8R1497R2Zwx4zNNZ3NUIM+hoWFDhK57d3LpCJPw1yW5plUD2TeKBQL+9TXMP8FMbIHnd/
LPAXz+YqgaZrOYndzfdRv+y/X09SUSaC9qjv9UqcL5z01zWutIGJkxnLU6SeBsvFdcXbZa1UGR7e
4L6rQl5GjPs4xiPj6MzJxhaJ7Zd4vnhgfXiKOxZUpmfMrnqiRfH7F7HarDaUp+z6XuMf6XxyHXct
/PVerrgzsZC/MqsKPtnuSgCyUZqrMsDJbIWSGagB1oUXr3mGGs2ZqhgQT39SbqoAr6XOh1SjT+vb
rnj9AH04yWld3rrhNUmyLzw7Iwvn0QhZCjvHedlYNRg6R+h1T61sXZXxbR+x/BI8p7ueII+aPexY
BTyZgwllMjGmsINoYAnGvywKGV5sld9R4IDZ2f3VkhS4D1dcUGwppKC0DmQ3y4m2ZNiTi63V0OVz
Z+WHWHkCtn4/ug0G8KLAzZDcGgFQXQ81K5FJ9v95/Nds7xQ/0e+EoX4ktrTGSWh6B5KMoWBF9UwU
ko0RC4r7kqo53voNObzGwchRa2YFWMMk3z+TEtTc/kuQGQsspmWHdwSWhdpMMMw1IPXXeBtJAQP/
4Pk2frpTC9a/nM6/baEFqcNqzk/eIqlWA31/54/wzuhQZN2xvbz0DT9oj23ACROPURgEDPGsNN76
TYpNTRvJtvMA69nnsBqWHA191d720evmRShAnxJM05v0xL/FMr5YYed0BFoo/TEgJ4emc4VkZelY
yWiMUciHTDUlrsT1W6HEq4o3zu7Iq3iRXY2Hputf2qbENO+//455gap3Tin+3V3gQFPsvbJY8Hz0
EoJm195QH2Mf4QXJOLWdz9wurbFyx4Wa7jhJiU6Jaixm0NM9p8hG+9wYfLnFmf5cclUsGBQT2hDi
up7SKN/xoRatGFNMo5c9XJJAwV0whwFC4d4s/0dyyjPp8aP8ZTQUDm/J0iBfEzZ65qRT3IxNsC8Z
nhzSBW+kwF/JaGPXBpkobRBKY4XBUCv46oyrTl93B33YunmU3kMUsaVwZFWYS/0ZcQuVw4xJTl1R
6SFBooUmrbApjTpQq8+0SL4khWr6Cn18rzVVRhWSDy5AdL0x54EPiiV+jT+oj4RPrhtr83aQyl5Z
VGXoxznTe57W0okchA1Nxd5AbRd9nFL7WHupubh8etZ/Q3LrzADP1Cp5DjgwWyI07pcuxZJ5hs4D
NuL1YqQwYsAr/2Ps6N6dwLBrslBMRpNsYqWb5rFIk2TXJ67UesOZAIeQJMz/7NFtSAOpjbELB/8T
A+TU673vYpFd9BlWy/HOSSIaJinPHwXV7T5qprexpvJOJwDzvkdxsU3vK1Jv0SndSh640aC4hLVm
waf1MoRjHJeWtzTUioK4GpegatXz99u5jl+8SI7xQlXM4N63soRmwt8jYAX6lj5HQiV8RXLkQiki
rsQKpm1cf+dRxyyVhqmRORgUlQTMWRxGE6Thb3FW1k9EP5XqBT2ljsMe6mJlPzyoxyOdpiGTv8Rs
ylOIf7x8Pf8WU7GJvr8E4959s8cm0bDyKA1NCcv6S40yQoocGmepq6GyrZCqS6mt0rK/pRgzNA6r
9gXY/QUA7mUf5NZR1BUii+1/nXsULVbj0rR2cFkJJFgVY82dokfe6DxI/NPr7S+TupOFYx+82ocb
oepp3X3I1EhaUSrSmgWdKArLl415vUmtqWLJqnY5g1hniHpSjJEIx1N6MvKryRsePXENJfrZ1AyJ
MJcObxZvt0XrWd6v3IBwcuBIAuwY5JgSakA+CODjmCazcIQdrW8JAI5FzRYG2yCMcheBCa4wo5zj
o7afudJ4YcIbAE6reVkoEK/dgz+dq7dIt+GBJC9q7/ULAx+qM+AkA4nh38DN35WOf0nLlaWEK36U
rcenloD/jLfg0+zvroPKzruAXA1pBxSS8wZI4DJkObD/xAguwbbV9pOEU7yzPddbGm8Kz92AHRF1
7kfYuVv9OLkXN5fJ2N1zTZzvbwHATApZcNthCwLXj5Ixo+R5+bE21/G1q3TpLarBe5YoI3GZ0m0t
v18YQvb4JXmWrAcusSxWRrWEp7OBh2gXGnI0P+Kf+JU1bBQNT2n6yHx78KjSzhPlrfDgDk36Vnxy
xWh4uX4gqqhPk7lgmf9FFfKoiHsS1toWhWjC4gPSlQlD+apHS02dOPkM66UEykxWCRqsaPXHknwJ
LIfvmDg08kugSdUBvcL0INnME5M1hPMmqNWhGch7vdPMLStqnRKoRaxqCiznaSUxeWCi+GRUxF9C
D1NKxXWFDX6dFJjxf2qCwMmhFsW/sW7lflRqTJMx9uFXASQhOg/mG5ANkyfDxLnnxSnd+9P5h2lO
COqKxBlb/pyPLAaM6jgV5dW4FcxAa7eEPbbjxta3LOZEayseEPJgPktconpQ7ymPdU0k07yZSZB5
9qqND4PESHfDtl/Yq0Us00s2f8f4P808MIIvjvg1B3/EMXOPJLgKtMrTKtEeJLy4t1JCTgYL3qq9
Of5tSPIINdMypIz/xJMdCHeBNO1Gfo935vjLCwOTAqohoH4zxT169olPaY698QHOnu+xnc2GXIVU
gt4Iq3xKCqojf5rzlDMpDfNyLoT8GWl60c/k7635PxUrp5Hf1Y1QlgppP1ONGY9QwPfaiwCBnkeB
HUxlDyxkQaIshQHGDI6UM0Ak5PFRQlkJPhle81ueZtEXrBGYNgYmIYKepFvn3vawJWJS7oaVIhGy
Zo2gEfteHL/N8Duenc+ERN5W8IcPlgo42XD5V72Tpj9U7DLDreSZ0EFwDqvirhcNZp49Od/MAZWZ
UDKstIqN/WAayuLLW6lu0Z9/1DFdq3bwRQhHXTRva4JisjsTd70qebwLQR8QVJ15Dk5CFNQKmjuG
5HoW1rHxHkOYvphYWVUnrEsAUDR6O6pITCIR2KC1/lK9pfDWulWwVsWAeEPjCrNWnG0EqYc9I4eo
0iruaG849Yi+oHW07mGN2miT6xPCEd/o6r8WvK3+kKbhRJADhmPpbnHp2XMDQ9Lxb9VjDbY9jGmN
e4f3GtLPKM/twIHVNYX3+UfWFXIXPffyTjmFf2DiaU+63wEVVVeGfiavwxrmmRHBCzxZlrUObVTd
B32TFhKCwCAJQz7u0gIAIlDV37wVSenuW6Y0xMjT1MB2t9h3SbQx2Q8145+5UOs/djRdcpIt9zBR
oFrSIdY5Afb+y/yZvdhSu6JxzruxWrdGpAt9Iy/aamLWdrkdz2yuw9W/53W0N9cXZKbK1W8e9PyL
3d48YZuxWYfRxblG0WX0BnOwhjyIkkJoswyPfIxAvkPPJFZCE3trWwrGhvdSJOnRwKMbcr/QON9l
V3mruvBuzMICzuciWyszwFzndddoQ23zs8jHp4t+l877Swm0ce9X66UAu8LZ3omqY0UxBbDt4prl
jgTV5VSselwQoqlPkIXzoWecNGUsSPlLhvKoDgtzkzrhekWB3aXmsqbanqTVfgNjssr0XhSxWGuD
2heSRCpDSv0jcV7cflb26e9rJIouBRzLWy9rlEpDa2W7/PFT5rp3P8zKRPmlGnj7f/NDT48xWIJP
xYmMHgoVp73fGhD0DOhstarvfUVqHojijNG1wETHT+bpYupyi+sdyHSUgrwGTaHYIghVOnV96WT9
MVEo7hu7y5eAveuGOe+rRlEAtRXA8weSZgZl23XrgxAD9yRFTvmURlanvUwPMB3EVAAHBDuWmJrs
qEAEKoHpQGk7k3BbWm+HikzvTXkRNojsj7XjzntTkWhM1MxiLyE7e9U3nWGckEsK4uRa2gxrkM0V
BOWM8zoPHamMBfGexbPPVNsV9DO4FXxKAFFQaNko6w2R9maklu3wOZQXlWxmaRAs0FDUCoLfnw29
cGXnpzd4JO513IhsMuyMtssmyNQKPkCykhk+1c7eU3zPE66AC3mr+IY0UKEj0jnKXEYWs/XWjsWU
zATzwo3lnQjL4JlWChupJyK7JTZ7WkDgRrZ+lSZ19e0ergaHXvt2feOBT4GLZY4bIlEOqwYKB/4W
MT48Bk09aazHOOt8+WWnMSmIZg7GikbYQPHqbYQska0usgzC+TM18j6C+iCMCuygjXReK0ILcgLH
1dFcdMUWtyNOQcPhOh6+L2QZQ2a3GBSJ19AajVyuA8r/8kgmwEFGXVHsB09TiUwtxTPW0Efg8zB5
lNRrfOdgR9begnmhaxLWbuwSdnaXkfWo8vcrVGq9EW7r3dTdwTw10RfYyuwN0AzvztnscpwNShqB
h4i0zlT8lno4v7SfkUjcEhjvzWrFL6AiN23uvw3Ibj5V1mSCxq8q+cevF4iwgSPWO2VvBO2g6ujG
Hzjn2yKzIOCLAqFkStQrMT49tYWbQk8Zd1RcQ9wRJ70TyY7joz2fLH+LhrQ53N5RDgf8sDDTxXjL
dCIJG+lcpQnfuBYHHOEHqSmTtr8oBwBrcf3js2QTygN4NnXjlJFaLS2z8QBufIjCm5U+nW8OU711
URNKVP1Mgo2t6vD1NK8SYBnuhYf8TxQ5Y4LHE5yp+K4TNTOSxRVSTowGkNC2eHtsmWjfw7qDfhA2
uYWIBjVh1QsL0ulBlSM6hJDI8ApgN2CHO1WSQgcXSx46C18cbjroMLMbnyINXhbdMpLobq/rkXTq
BLbOv2Ar1J2fLsxra4O+h4KYK75dtfVrhoJ2BttEaprJAkzFY/v36KYSQWYhtPSdo/5njtrr6MMH
UuOaB+Ku28pmd5Fa+IZ0+Z9SR9rv4vIS4nXXq0H6YDHrYrhZoAGK61VotgkcYQsbs0FO7WB/wRSu
uS7T/iCPEL3wgDsFfKU33cW9rGAOMKuZyxsoynt9SUYoyYlUmjV/dnh6DWjHI/59u3jwIHE0/3Ip
F8gV4MCeO+uyY5H5rmfLuikt/IXajt2mdN1ullR5hbDh/QxsUtbPvoE9JGgbw3djFUsA83rGQbum
NoTRdN1XoWcNvDqQLfruSrJgIrPpE5rEtjE31d7FJR/YyQLCgXK6a8POCHBbfG2Wk9+rL+5Xq5kB
sqWc9CyalTuHvJbqAFtI7+bz139wIvZRo87Acv4rPAL3jNGJsHY4xPuKNrY3ZQ2ggWwDJZZKhQ03
6ql44cE+Gs6gGBfNE+bxhqnGKgaia3m0vjy9kfDEyDCxDYs+Rg99rOq8Qwhh7ecMjidcN4qSgf0P
P9/HBCd3vt5Qcj8wADFRpu4BWuv3LJnrBy498GDwWsrgqBUl8wU5GCQWFsjb94Q1Fb/URM1+2MSa
ZnAZP3dc/vTd/nP6z9AgdJAMcF80/5DN/4GSQx7FiKW/NunwcDWlIvmrfrKo+yvI1tbuUYBeSW1G
mQhh64kU6lUUpR5o2upx4Tb3TkjRi79ZmXzXBvvZwOXDMxGBlSp8TA4RyEOpcAayb/N0pRcJlpn+
da4KsUweDXrQ7tWuFtL1gVjJH8kKNThD3sxPvbRvq0u/f+tcX42gs32zxlnzj+sbeZqfTFqFyKMy
2ctgmawGQ1NbiJ0OZhvOwbSaqRG6mwz8g/Qod1nzlysM65MINnrGl7hCYPAgtF9Ui8Ho2YA3xAJJ
Cut8qQu9/agrJarOGArNLjNIwkSP5vvlJRRe3FHp4/MP7QU915SU+rVXufhCIMo/A0aGH1ujMX7P
o70LMHpc03BXEvErD70QjdvzbxyUJpOw7D30cye3+COkMnwwHd5Llr7Pcld83YqSRvhvpYxVO1zp
8NmctXxHr9Qn9wO/Vd/9POMWKjS6m/gZBoXrJGo4ps2VRHBWG2DHic93B8dIdXmZQQ7zln0k7Fv5
m4CO+U7C1CTsx9tK3A08/pIKEQoDrXE6GWUpRJIjOk0HADGo/z0ZsB53ZOHYc6yr+8YBkXgVO6v5
ctBeb5jFZ+U5zlRlaf3bF9ieq8FGTU8PYpXQr7K0bdY5HLcHsZY7oLcqx/bVpzUiTd4sUrjj3ozX
i+MLPRJ3A3qzsahgPFJ29uAD80ZEQ5yjZzeNmYyW2ddqInRix2AKfxOODgKXGOgMVpG193r9uN+8
pQEk9++d+Js/zaD9Q9YW9M+Gwd9bEQAm9J1ihObLMX67UwjBJRKIgGH8SLDSUeLmFO0yJ8rh1spf
TLwoZZtvgeBXedyMO48c3+QaLedk2MElvcVlWao+hYhmIwf51LrVShX00pgGjNDFnD6ajXZZaOcq
BjTAogAzQRwEI05P80kMXTb3K13QRpVIJGHrOoDt7rv8BOq2t/FNi/e9jTy9QNJhNKHjJ0VKbeZf
FJ52LtCkWyWJNoZzc38bNL98ztukvEA/NOKqX/VjgYLj1rLJGf6I5MCg/OTEBCEpf0xfGWrFf17g
fv6DE1ZpjvvzsA6aW599VlU1NwmFHuLy32lhRmRWN7+6qRNHakRUFP9Vjchy75FRLLwqOj1zAoF8
GCJlXam9DEpgwlppwbDm2uzywCHnrxRukX6sY+Trxq1onLs3ehXdeaWaAwUFmPT7vpODQcVOrR35
qjSRkwH9weMDayZnsLVh15ocK8iIHMaeSTQea4uYNuB9xcghh9dna468gOdPPKQIkNMJLISPHtMr
1IkMp5sC0yTU4O5lMogHilE03MJs5LajHmmTh1ErDHT4kbwO5rDJxxaFNX2g1Y3KgoWrPAqYYK2Z
9t3bG7Nqgyv7m0Hdo8Aa2sSRtlkt4M6PoxBk8l9gwY8Vzu/tmA8Jd1UCAU2+WFadsG0NjNIaCQcf
Yw+imLRqrsi0F+G54LtT1dFRsX8bPaZVuUK6fx4hwF8miDspMxbsFwNtD94Aa4AB0MSgNkcN0er3
KesJuERP3H3sz837lcD/XzbVODF+Jzg+UqJKh68UbbJPMF3dw+97qjRmxxS8aCLbssbIDjIt1ISD
OZFZdFqDWRxJn0iaHPSnBYxZTcG1EwjQu6lkB7JulTgiV8hGWkHJ3R8/e7cBEUHDgV3KIr5jh0sv
tLcXnrzT94aeQyj3cSDLZ6gj0P8RWuE4H2DktvBQLZc81G4KrCJpYtoVeqjzcAA/b6O0UDNrXjY/
XhKQEK6OVMPmuBx5enpaJ06iIvPJqCK9GTtoLhIKH71pxMJlYECSRphLDJh8q7gpmo1DrUoqWJ0E
KLFDHYI2G21qDoO3Z08r7DfkybBjSGMe32/NHGALfvUFxsrJMY/pq3sbgWmC+2AsU5/JYGJgQFXt
UoagAb4q/ApqPZtNajfRgFwRZbNsyhlpdVXsLjn1lsZX3gfhUzzSQs3Oz3zDuJVxIAYtGQZwP9sd
X2djEwDPllAqwj5vlB8aRvggSS6ioBwXd0SPMV+cfukD9NnFEaG+Kc6lenZxsm/d/b2vN5sHLiMo
M/t3U7pqLaG8bkceHnj8EngqetOsL+ynVBLfX6dIo4OyUU/3vacCGo1bkz699zPKXo/vGFhT/BCC
26MAOdA13nbq9BsdLEXifTDmHdLnMmbdi0H/ctgS9mR+0vyko520zwnMV+ycKTY/xzTP4O/BVUII
57pyW8lk1h84xrizhS/9P2C4RGTjtT6ia2T8nMRVADObG2N8pEwCQvDGdn+U5uxNZyolqCi9tCbh
45WNRWaZ2xKOof0P/pHmAspwkExCSt4BNmxv6XgKDT+HCHlAerO4VNTl8SC7+//m6ZZi8bktVhH2
LU6pV1tZWogYL6fN0Z/S1I17vH+90iUQxkJ3YBFU6WJK77uHDueOKc3OaSIVhAZj8OdHoVV3er96
owAKX4Hd4jW0fOvDLDYqY98GjCjuCWMlrzboufIJUAQYB4Ls2XUAU+H+xhylGRkF6PQSTpjkDoz/
DdQDrmsDxeicjWdkLmcI/Ls5T/xqbCD0d6khVmRpaC4Oewx4H0pDF5J6ljys4taRf7czHInWb7dR
k3Ax0URjJYgjQGYUXwtklTw2REMEKpg2kTk3aBJaqI53sRxlx6eiyDjgdY5SznLzptKZ1butV9vj
A/NFyp5iWWaLJH6ON7Jrly7w+hAkA43Fy1RFGiDjLAbUURLVCUVyL582A81UKdLqaqh0ppE/OP3V
9XIYJH7xy00VWkAgtT7J3PvYxkfB2ilsXDHlivEBXVV8vEByu8cSJm30DJ1E5I01K96FmAiq6YVe
f+C3VjS50Wrik7PNTWNYYNcVbf6Ryu3UMcVGJqhCU5SN5O65cEexU4DJsujREm5Wm9gzKoPjIsJo
Uurm7nmlWAwN3cN7OKWmzlcACfNmApWwqfnv72K1pX+DjDKjTawBr+cTHakIBy+VlUwjtYOGzDxB
M19AWyW+Phz2wKPsZy8336a8qlQzdBj7HgyKw4Ptbp2Bzx7xnnODuNXE/Yei7PMgQ7wXt367yCv0
MygfsEpNFy/cDk80dZ+AamS9rzabiJFaPPYavaq3+Q9eMiRKEhhdS3sHLuT7pUhvH1iuhku1YLJd
ySwfJgw9xadjbL0uaagy7tI4YhHceBgBnQR3+2+LFXWemiEZB692we+WFG4I/PPopb4LSRT/uvPT
booKKNjOgqWwg5B/0w+qL/oMCvHfKOz9zfXIroV22cyHGucv/Cj4yYuqL7tuTpl6YsaGdKG0z7kT
BhnPEhRWTebk3/RF/s3dZphu+PQSlIC6uWc8wXMPFB5B/0blN33rI2ABGSGUJ1ndjE9+SoL8zUrs
rtKxhKcx20yZ49t4LF2L+AzbL9U1mRlQ2qSKBN8Ze6iOZRgtMhMnBgztXRVER1cE1qJnQIqnxUyX
HlrwmlIzzLgD//qk3avNG977umrMMuY56IH+A37mAK6a7ePmSSRksh16uUstYcLo/PNwKp3W4Y5h
soTme6OM3tlCkyxnO0/gT0JMABKcNDos1vFNpw0opWScljfmsTq++VnQXIcvnUZxqdw8esAKkeZk
ECtjOgQtKc4spoEq1mAXyB9OioKY95QGIfXzvLP3fKhiIg+v71/dTAid8w436fXEElyjKrijpqEc
LHrLcw6k3RO1eQpHkPv5xEwJ5A82f1Lmt+EIzSOVf/Gb0+yM3y9FxS18LSi3vPceSsx4Wz9zOVw1
6bmUWzwjQG0BF9b2TtvSiUC/sX2RR9upf+IE87kU2ckLYjjvvratDzTYkJglrIKGzqzIMoNroraA
cTkPyvDdb3hqh+G5TquqNve+8Gkr+chSInk3bAQFI/gAKPatIsy/nofD/9bx7g89g8S5E7ss4nXz
VwSrYXYuZZ57uhTjmoYFu91K7f0Fp19tmMfWFhYQ92yt6vETpfgJ8KAgn/xR6FUrLAGeJ4i7oF9s
/FEgf0pUk/oTyE3R8Zqk+zR4vImtu5uagmGZy6SMARdxSXYVJwpgLgdeahtRQ0adZd0LQNALEgR5
ZZahl2lx7bWzG5Pl7xbjTYLol9fhocLxMX+w5Zj5h8wsUXC5FLgWDCv4G2t9D6jq1kQ0/BrF8A25
E5Q+gWQ5tOUUFO6OENtv1N8OWCR0/xpiyPge0r/hxJeIhTMtsEhYPgk/b5gjYP4ASku3zpMK1hTx
EPhsEOOaLhmyGylXVa/L6LP5u81Z8rMggh4JTBBI4sUKHF7K/ujkjVT7+S1mBIUjVzQs040EDK6N
u7/E8xYt/kFqHaxsK7ejJZpFvEzeJQGpVOGp8frShbhkyR7JZIH4SHGtDudFw5UmE7tjpA7YGsfC
q0yM+sCdlL6fJiq9Vg9v0Wfw3pUnfB9X2Ak0CBQOqXnBnxtkeaO7UialH/3isvMJfC6kHHhBTBYW
BL8q4iZpQC5N3YSG17bNdUudUNM742tMSjNCoy0ecBQMuwZADr3M6A/J1M9CBM8gUhgiJoHIWr5i
S/Fb2dUEDSBVdIa52YvgiLcmOfF7yee1LlNMkVt2cfgymrlW+xfR/5aJqE5mbh3HTY9IlU3xjKrZ
qRiOwG9p/b3zHOVqbTF0FnVLkiOh7LrIPQOM2dMwf+Bj0OpgUa1WUm7vd8fMjkvwE6VQP8ta6HI3
q3sgtDxbqUF90KKLwkz1f42Skjoa+1vH3ZYMuZ/ozmTxltIjMfig9wsy/mbJNqzYt3TKCJLXze+s
dMbRl/qNC8H+M9+96yDbxgnF1nzII1hbD1w2JgVxcdiOXWydjDJ2OSjACUChPwBzRVhEQ1WcNe1k
5YTiksv1Bb1efLV4B7wAGtZG3w0dKcPYhCvL1flU/ADP3EUH2lh3iEiF9RJ4lD44nTjOzuW7375i
l7A9CEzhdnBRln2NxB2pmsnhSC3rgDhU98UJ6sUUm9AinSQPvCYmTJBCNhpXedOEuOsZTqYN+IiL
rCb284SGgyZZ+TTIS84sZmopKB90iDJqWuch0zaZY57jcclijvEHwSmAws6a7c6rAn528Xq0dk0/
rbtWtr8mIPp/tmrC2cVB5dQdzyyvd3M1Dy8/NxZ6W/+6z42W2j2PolpGTYF23e5HcDZ38SThf7Zs
J/Pr2FBmIpcD2QArLHnsrAi+aUNCjgaxz+ylVn84PL+K7mXSc3n7YiyN9ZR2vY8U1Q9XW5krgmSl
eqQ7p3OwMbYPfy4HlDCkHiGEK8V3NjtTSQh5Bit04s5NL9/kg/uF7ka08HDEcC4YfqSzackZt1xe
UcY+e+1x4L/XdskwAYTNL0StsYaRPK1cot+XxYyIULJlPxfu50kQndRDio48AdF0E53QcETQjpy7
Udi7SuoLfStdfXMQ/rA2uEkn7Q8zWv4GdVSFCsyQN+fbTbt1XEdEnbZlBUXUouwpDmKIJ6oJyIKl
sjT+cNjYru2WRRw2pC+/Weqm8awWlr/nOGNgR2ejZRKOLc8jIzf+6nicNDLaMk97kpI2Vy5km9sE
aKsidYD8cRJfe7FoYjs4u7MxbMCLmG5L+ErWe4NuQWt3AGQW0sEidDlUklOzSlDjOw3TGXMYYz6V
qKE7XxyK1hZMkALXfjuqqTN+rp3M9ifyMbhLerNMpv0ZAwhtjWRUUxrjiorf78Yr4aUDocTGiaHE
vEL3Fa3Q+NnysfUsDZP7XZbTx7Aq55QrxrIOtvoiyrrtP1DUgnLmWeuhqUDBjt+QqvWpdgNj5Q4y
4mfn5awOewannW+ln4sARRLuHfmDTpS/jkgUgpGm2nkeh5MDfOIBS7qihTQM5aqzWnaF3bRwTwaj
ebMf/LUwAwOlDAkQrR0i4tm4J+G5YdOReIL2axW89ec5NesyujlnMGSuaqBvdZaozTNzqf/z6cTl
LqVcX1CZmraVtAMW7qSlqzZ+XHBYi6/TTQm8/pbOWFMHDkh3OLvtTBqhw+FZwl4OGtsIc/TX0X07
co4/mm6bHqjYk7VlPCmouidCkMQYw9NSjMaDhhtWGGZ0cM2pyb4t+1+AwgoqGfAchLCzqv9hZ8Ur
FyZTG31UT2BptfgnOmpBdR7E8pspZ91U14OKn8QAEHoJBpn8y7BABnpwP+K/DG8AJBxrf9jMXpjb
+K3ySmjG3rZ0wbqFmyfYInYkpl8JRevK0Lpgse65HPL7Zj8mk2ikYUeiVWxCeEsarw9kru5o25iL
g+Whgt0RXj6bM9L/Jbe/VKYKJJMxlapqK3Dlzsp8Ks9efBNmKSZqS5UaZUuQq29v6IHyug1t0LOB
7QuYcnmIQh0SkFQFiRNwwvBCxCtKDQeI2zCwwx+Y7OvMFYblfB0EdJNESDDQdRqCdgwuRU+kADMl
XFQfYH//6xDYHH4K9DQ5Vyd9vNS2iCT4O4pVS7VO/Y7d3wtmyq5sDs1JVyMWl2o0FwoIfNUgA0DE
auLlawjAiE+zxVKg6i2zetTnZrXB2U2S9Mb4JIikKb2aBipDZo5IIEPCPniYX0jjA4NYmMhHHMZ3
flPuS0t21l02Oq2sbR8m0MDU1Fgj3VvtXK5a3cC6J9O797IIWD3+5UVdPVHrsTYKZTS7zf4GGG3S
bmplngfrDIY2SilJmE0NgsyCZ/w9mfGJeeF20XeEVxvvRWLqf1eljeH1InsO5pxN1rrXC+pOtf9T
whbXP4zqa47vXpPdQ3kQlJNGv7AvlfZKNJsovFZlohCeRpe83i1us3YrHHGtZSE2wVUU5hFFHkm7
09mlPzIUENZNKQKDcHvcyvqq7FejZOeC/4vauHARycrQ8e8gFmSARs8B/p3qKfFF7nyAp9o87RVZ
2FkZLibMkb1g9ZztMNF1iz3K4pKtwP+CQ/QOueoAuhDp32N+T0si1ENHFXJlu56x13TxkS6iRp2O
MX/Ec0Ff5751yHE/VpLMsXrXJ/KQLmYOteWYnDUvak1EO+nxvt/GvLFw+GHtOOQebUWW8wrlCFt/
1/e63fhiQyrhH8u2WZelzpQur8CEI/cvXJE5L2bYtBw0juSlQeON64Onm3n3ocXC3DVHfNXDa0zk
SB80YxuSjEya5W2AC/ZkryY0JTLoDEKpaP+7TA5le0UkR/smsoJJmpoUBMYAniaFCAQGnhf7uTBQ
AUGuhd1+10oI0li2cCNA+fZWFGtgAy6Y+njvKbHgydd5HHFT/A36YYyUuwsxNTpDwoAMbuRvyZve
nst3s/T9+rKBw2xL7N4SSdT6a4Qe1P44kemX+yINnx8rEbcZBmx9vjO2bar5Lr7NQujHRcF7C2u3
09an1KilPB8L9mWfR0jrMUOVhzDqgpxom8pi3BmOZ6kTogNUjwDGps0ZyATB55NzpyzMwD7JkfWk
lLRnkuRGzTuOBK+lcq25KxikZzLpzK3XBKWQvBbwQLGBiTh0mgM7OTUZkuOUJceVWQGMxMFvrDDQ
h13qcoKqJjYn5Ka5T/M9VSNUO7wq/Y5THtUxOVY6Q9n4V5c+9N/NVEud1xO5F+/vyE6l0wXZp+w1
4fQh8/LdKx33/TV91hL9RSa1CdLge4DRrikcLlHRonXWrqNcZBkJnAUekJf3xppnVTwmAIgUokZz
YkpG6MIn4dO/jFEAjkR3siY9o1FpZB2TslLRKOo7W/gpQ5LvW0K33NytcWGoLQ8+JWEZntnc8o9X
kluuzs5Cp06cUY8wqHk+3r9YkjmkTWpiRaLx9YiOOuSiPbKIbfrH2lGomfXhVTO58uVdA2w0ZZWN
WqB1FD7llO9acjg2LkTdQVm97+gs/DtQSKmlEaP4XHoGmt3D5Ny6NJzNn7NhIPjxxr0pup/w4Jwx
FRB2ddsaLzjthn0sG8qnoz6AfSs9OvcAj1UEcsFQqt/VKENIDS51yEW32K/n4eN4/FLY4mDMU78o
RRoq8WlfTtc05AESYGuuLPo/Vb5gESjB0AtO9rWQtiTbIL2/zDX+wqWiaYO217Gy4KqOMSZXuKGI
vAvB6yqJ2d7X+OyHuSJbRQP5qHztgMWdgpB+O1L0EaW/YW4Ub24JMvYe7t0xTYpFNLDya8CVdgWh
6Wr6xeP5IHkNgMHeqK95tvCCJQ43d359vRTEfEI28lguuHizgsVQwFRCEljOd9jzmDJ0Y0NdmR2j
jJ1cZ82dtSKr1PjU50uqOkBb2dB8SNiJW8d51fWJ6tWu0U9rUNcKzAQkGUxP1hPVjiDIMx0bI7wg
fRlhrtkcoiOlZotWyS90APIEzrdA2vieAarCosTWJvNAIYputGK4/l2Xxrumx3VzxoABGixYrxbp
+YXf6GvJgmDAzV/s3X+j0nju1hXyXtknVN5H4/D2VCWjyGUpwKvcxBB0CRSaqtMlWkE7hUVoiHH3
tDe1Tp0D53PqOquOmOn/34YDxV4uAof4m4YEYaZpETo0F3CNKxzFUD8g4MxkOVzXyqofTeahoIP+
7C83dFAwkX4enImehab+qzO6q7mCWH147v7nTB3wCba/JouN/Js5uXDed6btusgMyuBOge5Wdsmm
cJE2TrRGlZVIywPi/Rb02GjiErUZGBVbGIA/RAwBfbr7QupCufo+5cEySdHBs3cYIoPCXB/SGhjb
K63f0U0kyTlISl0lTZK/94cLLoDl403egClAs6ejWEeNZs31trCcB8v8PrhB5nOYEdIXNYiKrFYr
XnRzZ6rHXNAJgzQDnYSj2OjSp+rqLSiWt+XpfD0yN8jPW1QajH1CUXqvjgzya78XSA9Ov8IVZQYC
fG9KtaB/hWC8vmiIOuuiCXU1rCWTrZ+R8lvqanC8fGERWWWk0/UCOdtM3O6NnM+KxHAcx02ULAdb
gIb2Ovv1MeQAFPXRM5hPIbFZXNFP4Um1nflV8H88QeHUsHEjfOoYqWE/whC+Wfl4wzKSmH7GKUSV
QukLryb+VkvDMh2ht7ubZKINpbIwpIOTne+oKmBka8bOAioJHBllONBglRsnGGbcy6edPeTyJeYk
kvnWjJFZmgOkJzfiOmjEw+y1KXkZ/84Mc4v8Dxc0C9MlqjNyGlYG/jl8j36xy9R9slAy2/NE4/hA
9G1zvvJVPd5md7Okhvgk8lrSVRRoyMC7qayKJL9psqkDnGqDz0MgzhZZz7bhdt1nCyCr/8xJNbqU
eNwROUGIRPFbBXoPOTOQiPH7tDqZuaUKBX5ar/Z9Pztiddl6U4KrpDT7Hn3c6CjDTC+E6d1ZsNa6
qEKVDmUvMytZw20kUCGMuWd51VyJFJE6X5WCd18vaKU/nhVUtBgnyy1InPcuThC41vKUCjeBoTBi
uImC08ZvpMnAgwabIKWv7pHgtRx+67lsmE6MKFaKw4Pq/Hj6pajlDEEfoau+29dvX+myTt+94OsP
HZSiiFPDrlzhtZFBCGlD2Uh/O86ruzEqsBPHcmh6Q1oN+zLpEJTpwV8V+IBOUmVehvk2Kyk9wRSg
pYl58rPzlO9EMjjuoeKwxYpjSdnT6C/6R1ZoMA4Yjzxo3lVlddCMFBdq6SpYcG027/gBK5Umo77x
n/N5fYT80m0HsafmLyCUjKfafFO5qQk1/h59qkbqZymAwRPtdT8wwGQHXZdUcLfdLJrCdkeO/lEY
4i+jNaC/GqFiqD/CRu3ggaKwYXeH3WtvUgeTLSrMyagBQojIwG33ZPDjZGGmmNAEfcrJ00p6a+Tw
SRD1P8PUQCJOBsomt7XboXAVFSNhGyKz6El9mFPfg7kN0igDckFUzFkHFXYV0MbRp7o9U4TkL8xq
kTlD7iCLrhVO3ZgriKzcC2AzRinij3F+j0/uRv2o1Qk7atgmz64OZ04bWM1eadqdBSAwjd5IjSsa
Mqsuo2pM8W1knaqh2IkoBj3gLUa7Nn2FGLuyU9wGhuQm4WyMrRGpMxFiaLDfe3ViJYNrCfgJIHac
/oVCBDH6Fi3P2jcnAsW+Cxk7ClLIs9PWASHXneBfIWvi6rtDWrTTbDGgPgHiOknh2xktEM9TQ4Tg
9ZrCXp9ZcsE73flF5H0HP1DCQPklrjED9E1cmvtiEP5K9RwJzOqmCyYOYSqcpGF43Agt1KUK2nmj
H+SP1HP7WEW3Lv30bKPK0KzDr08eVAwp0Ww3WCSVL1eSbWdbu2Vpd29Nsjx6uT1JGNBuaYEv4b/N
h0pUijCB8E6tnGOiaWxnFITOr3XuYDyB0hjqNGHKbS5rrFzX+2WZbSB3BwvUTuu6kp8Dyle9fGuE
iMX2K7qCo6ssUIGnIPofFQE1BFCpkV9gLo8MzH0UzvXt8bbvQyc1HEatA46FMH4DfWLy+RRfLWUJ
4V8UjvczXly+NrgCZVsY+2T8sSBNytO/0CMz6Wt8BPJUzyNlHyD3+5aIAjokRqlHZexfVf+X6OZK
zvH3Yi/uDWHJsfiLWTsX3qa3xN7u50LEqK9Fj8Uy0VrEyM4lyMyVuZt3ex0WZtah21V7xez/U39f
yepBQWiBm3mQcvsu2W++HvVVMkhuFViWp1SFhwFkhtBpVobTwBTZvx/K555xn1Pa2Du0VbZ/ptBD
tS+/Q5JO2q6l2Ep5RsvZ2Tn7DK2nVwm59RsbdyNvBezSXuUIZs4xirNfVIo49a97V8MFgFT6mMc/
PWBGHskp2t5KFa1/ROuzlFObT/lKblruMSRxxtSoZs5WxqnOrKEPCO8bBYlhduZsf+5LI4bM9XZw
/NB+0Kyy7EXTaPfYMP/HmDDKDmvOXjpfkiMJbyVJtrNftubCFjxaIPviRKsyZZrA5AOEH5hkpSHZ
KO8FOy9sLH3tKJ36wSuRDgHQjwK6hs6t0ZgStoqnv3nUFLIgjZ5i8s5rLv+rXOS8ji7NSdeX9vfD
rAzxyS3Ci53PcYaOBIKRYiXmf5fjJ1OEWph7fTmo67OokDnSxPxf9VqDpjoRWjY5e1xfwVX8gEBa
9YBBE1svG/QKQsIaH7N0Vo/kWDlCMPY+ZEDJ5RVkNb4iXTqQW+f2wUNJEA3wXB4Q3zMSH4ebpoBQ
YsgjU/OIR4FsOFcg6dlDfEXPLg8Ix37fuBwBzC8M/BZMDN/h1Rrcf/bI+3FOFxkdnkzjGoTfZjaG
opa0nKyqbDVVBuMVIyj+y2Ryd/mPz+CZXCsyn7UMOPKxaI9cSlL+zDifMnsxr7EoVYTantchRk6C
78TavSLcGXKdzgyHwHcZ9+/NsLlAX8gMI5oUsxx42VjD4rX76feURLM4kbUiDTLAUgoN+ISyPaJP
fhTD9am1AxxeN/vrzcy7JhLiNwsV41fcPyVCIFj4tqodBaGLtZm2by64n77KklBjTladMNM2Db0h
95J3b87wPcARVwpwyMw6EPOqRzCkjQ3k848RCxO2cBo6L8Vy2udFDlDGZnXzRwoQguhPlUkBidie
Pl1OVYyew9dCbI8aMS8CVpaiULdrp0ein/trfXhR1hPNzsW3tvk1c71tKEgeMi5Nuhrz09/PW2ZB
ZRS6MdmdDftR+klz2l3DYLY/8ExYH4jcH0kWOhTrBoIPhGMlJ884CxtV3Uorbkh0pAGT5XEzDPkD
J2uwHDYYSEktZ8WglJ4y/OG6E8EwNnDOju00Cc0Tww58Dav7XTF+/nGm98XU/oeqQbpjh8lNDail
tet5AoKBeicTjB22F1+LOj+w3XNXkEznNXPpFKtBirkVV1EOzUAvVjIaZk/A0N2uXQqKKedvGx99
DGA+ksv7kQLXuOnd+m+1+ZysoDgcVXgICj9i069a2ncZ/cE/PL25vUeEli5im9ITasArVxb/B/0d
09FmlvBJmK35pdvTU5a1n/VeIMLryw7ZfESzEDAyanSL9+eBU6EYjg1Ak3C37JZvyK6sp6UDbOF8
FUPZ4ls4E7zS7jv6lotJgI/iNtOd6wDshkOTMr+W+fWrMO+TQiKCrwaug0CIpwH3GpGOPCnfZZjs
HnnUdFqJKAV/EBqEdvKsWQfViSPx2UQV4F5gDMTJpXiSat77RGAFayMbmXAmdAUCIk5fBYe+/znh
9kuuvRJ861faeFWPmuq4r2eMHGPDJtTV7W8bIC4pUPMFJPV384J+hqMvkrh9Wzyn6P6G6Wks/B39
Q1aMVLfIelNNU3SskbfOXrnRz3NZG5Y5TccTm6bvX4BHFZkQrzav5T5ecCf6qeTAis5SKws0sCnD
NB6VmOpMXjC/marI2qiVkZNVPIymaKbyaPfJqd+V92KbAxjQHTeruCiKlTd/X77INS+PJhAheIg5
wAVQkJQc/yw0CO5oqnqjQdWWaUKZqhk1pQkwjbUT77BmHN7b2ZoDpb+KNyHrIs4GhDTLiS0Irtzh
ByfnSkrenz7JFOZ3WhKtqWf/otsqsG+5Gtxufe9rK3An9rilPrGYVXx2aVx4TigPzai20kbe+L+x
RwljmpcCTVF56O478yxYRXAAgCukI9qcHQPFWLR33LD8KUC5yCkukunM7g44VUIeDmTffKA0c4zU
NTmRP6miI6xZluWa/WT+SOVEMI1wH+hjvgKhjSxQHxk3RH4GpGviQBypjDxRTyrro46oUSnONmnA
ZEeC/vDqVRfGrUg5/+Xq4kuQ8FK7koxtxAVaw7nmMke2vw7PkjXZmV9h7xnKbtDwsDL97mKJGz6n
ne5p7YgQqPxKsswvh42Xh0XU1YmdqivDopveUR2gkRZkV0vqtMza2aJ7bAK9VvIj/xJJfFfiQ3Eq
K9IGmTdhutT2oOkrzh1yqG49fFWGSWoQHcB/8/jx1wr/gp9ZTa7GqhDv83A7BpbO7AINZ19p3Onr
DalACfjWkHj3QwqUx/VbWu1q/5MdNHtj16+zuAucjBreAlguVRQOaUguXoUVboBPrFakw+2hGURu
NmrXF2z7FeTneIApF6M+SC1Xd1xZo3ghMnDDoTpRca+gl7SSX7a13JlvMwENzsy/B9io3u/gzCJ5
DMzrtMxlt6Wp4JGlpSitNxsnFjXF2o8/QeZ4KxCxOjjcqjDgC9DioPRIRWQZb9KJdfRNEmEmrOwd
B7UWOVx8JMcnt4sM0ya0V/L0i+Xizc0Fpr643PPLavSNrWQZHyn4N0goauePCfXaIgaGmeSvaapC
KoRGZE0P8N0XnqnN4hnxbbCe4eJK96O8fr2mDSChB1IVrDbhiQtpVv7ndK3UmvuIzpnntLRwEBls
KdeTftz3IaBl6bF5HFt7IOOfErQhpZGTE05dfVeK5hZVQcIQG44sLSKMEH9dWIFXaA1VB+unCOqY
MTRhc1N3sFog4+5WMMja9Rry/Qu/RQllm87Qc1m/kIZyGATpVBdgaS6whiev3DnD0HW+9vAtM7or
Jbou/m0iL7fb82qEN1iSBMLfY/y7kXjt1icSdLygzzht4PID9HBFQ0b5uFkFQGCF6cge5WiimNLb
Tki1+YBF1x2Q60EFPkOPRZGzqjqY9YEzjfKh3zfDJrwdT77AKet93G5cTvIMrMkysZQbMweTSo9M
y4YGOFT/shv3jMV2TW7yTeKNUhA/stf9iCK2HERrGSxOBlbI1VTV4klVvC2hVDRfNkg0IEuZ95+Q
byQuSObe2bNQhU5NNWr5WHQ+DhF1dNyMyu494rCskXeGK6C2/1hycFeOCBS1oqDA1/nYN9cWnD4J
z2cOUxjaqGedxPYYFKUui2nN156RP1oy0/HO08J0fixWx2dpDQJq6SCVWn9srmr/dkDvyr5ztnFx
L4dM9ML0BU2q3PsuqTZTvG6Fu0sUNEuzXPCt0nHre82LQRpsbyvqEJ831p/858jNsfpA25rzKuaf
YDPDby2g/q+eoLJJj1ZxYBv1uNK+n+17J9LTnpqrtuquSgJ/KM9X1iZLA2JZA2avpjUnmGJLe/05
uBJU38RdMYdrxKYujXe7xX4azCucQwgu3NM1zPQ+8IEGcD5briCKaF2IPxxGqZ8MpE5CfkuQrG7o
OPHo6u3R4zIW3B3IxMQ7JMoanKMHDih0og2S7UgMoOcFVQLO+9WfcGO8uKCmxWtk+rz3WCcvSyyg
WDd28U5kvJKGtyhK7LITLO6mJaQk1MpWMEUg9emyJgfaeBoInBM4+O0KVNBGTSTvKi+vZ3f2IuCL
5GY+2pwbIMQOV0Vd7Sd8kz/Jxc+veM59o+zkLWV7U3+2FBumH70zxTyWuZx7m7+KQbFkKC9W3vj6
RhMRtqGYOCT+KnXwbpzoj1GgSCP6mk8Zczc+2zQOSBUYhScrDvUmZzlR4S0QR1vcBNK+EBXa+Kw7
EdumNNkDLmX4ivC/mQD1oO2i6PfboOZ0Ogv/KmcWafDW9YlwVCx9aSGCbXw1ulLrDrAo9xnJnXEb
XXvIRCkbqwsOgcbbx/TtC9l4SdGqytjVCY01Wc5ryKAApE3I12dHXIQ11wtScyO+ohom4M9V9Mbc
rG0h/LUXTJwnDFY2UnrDrpWRlO7rbX+DuzLpGjYVSkE5iqXq81ED+ckXM0VbaDSesc2/rz+M/vrg
qVMqqKhsInVn9/w4CrdrihKm7Ww9aCIAqygyQfZyZr8QKFlcwJ5M3kXh07MGA0wVreIntQPBh0JM
QcJpiV7Wc1k11urifdg5xVEtVLxTA4L53mVgM0+qp7KD+NE4VrE5oCeDn3Fb6hqAWU3+z261xAaK
BNJJz/KY+3JJ+rMl3+yfvg3UgyvMiWdFzzWs4Nu3ne+/Op/J4ggwAyGwY3iG3ufvVArXtOz0KDt7
Clifc5WIHhGKcZKB+p+Hi2vLREI/Epzif/0FbyoA271nXb5CoqAE+Kpqo6VC/b8Mba0NEhMkTZD2
t2523oTZGRf1d3UkSvXkBtzmFtLxV/1Y7GalEUeb8XCMPjvkmRcHZuKgWebGjsOAZ2xd4M+KfOSt
JKNerW8V3MwEdLPJG7PhLUMuniYnVS4XWb43mpok+ExtDm6wt7SOXOwuMg0Hd5fEfJjbuYgzuNN+
s8an3bG00Lio24ubbzRaw4fskAKwzTATWW0fsqYkW2YXeq1DvQS/J91DLtAo4c4hwOFu1AwXR5/p
oMwdh5KwK4GsEBmDBuqv7FpLjlcdHrbHEalPRbDjT6tqqKpB3OJIaZpYjE81RKighcNGXIt6qKOX
SPflRPW0PKPtTtaVWA7J6u5QBueXTh0+1BDe+BJalefhmMohlo0bCa6iZglJB1J9BmyDGMSRsJ5N
PKscOdk5Kt7+OGhUe+JcDAfVsZ73eSUnyvdqumQvvnqdXlH6cAwdz0EDexzN/RQIxObiDKV59774
ho12+JMa1kMHo05/evy1rbWt8y7Jzd9dvJ1Q5vnmMWtuEoQ08Gt1LcWqTL3MtBZeKworHUZXOHs5
VDnpvvtbMaLKX3z2ymGysSgPcKIw4BKa4WwSlSyoWHAlmTRpRJDb5LnKsO3+yDONqGl2bQk3byf6
hKieg8KYYDqrdeHdLoQufJ0Icz+I8UZcx7AQOlZsN0c1ALTceE0Fd2AjygIjpJOHpIJPDmwC5D9B
6W83FIS/S/H3p7BcOycxoPxf5GUTBq4OUXP8TnJIVqDBwexra0p7/ugoFaUc+BiCVY+V4U+htc+d
XLoNrnkS9/8yk1Rw/E11f7yXi4THKNE6Wg5hgbPgxLfdIo5RQC2G7/vOa+UVfcFON6HAeVRdZym0
ZG4klS1pXLn4GQZdbtK+c/2Rp91PBoz2PIMaA5S5G/7wqN5e6VqUDv4fgCgf4wSiBCLJU4HYLS9Q
/4HK/6eCr2xhZnIOo76lRWeYUYF7cprVZjNXh1LlDAchtXZ0pXKlJ1og7bXaDUcrDLZU/JiA9iBC
RegGjnohbYxZySulV2Goydr/Mr7OZRNarD1yPORSuPB0FdzTaKQCkNQOThC/X0K5ohihtivWG6nN
N1bj6cUpi0xH7Jons0nlLfY81heRGhlrkFEgNkOlFTKpCTurvxU1lTc7i8q2F2CS/NllfitZylvC
Ft2VHEXzoROPICtoRH8hqfcCPlizBnwehQ+Req7WJqVtU/KBi/lWNo37n1oQyxGLY5Tln3+YotB3
51rFO77c334NL+4BP4A39TN5mNDZbejQW4XeMhVhtJ5ulplZGOBAwQXXE7ZPA1J0dwu4YyAj/FwJ
CHazCNqhOKbkxKeQbUzBSVWSzH14eMP4LGTW4OswNUQwCWLJTJkqYuhbaw6jiGNsNiAsVdOT75wQ
BrNTHpQF8+V2UDuANzXkl0C6eSxrzk1CqQxzKD3YijQqV4t24WYNht1RuAdZk5Cxx0w7cJAO3G3h
bfSqX9EhRL8ZyAMDDNh6zKvZsUN4jlWnIhiHGexbCfW3nf9iX9nMbnZ8312fir+U7BmvcMDUpi9A
gIz7ArHLejH5FfGEdLTMwDBafVyGX4pi8qDr4JFOW56K3WkYuTYoazbaoMOsKx/w1ovruEj5hS1o
kVtunKO3B8p1RAFUztXStlqUc40Ytx4IsCsAYPOfIbP5Hd+xnbQLy5G4HnskxA5i8KWoJ4gkQzVj
vk/WBH6EaA/5oIvYxbJPOY/XY4mgKRN5Cd2xyO6laCHYSo5QCrZbltb8N7npDeO3LozlqSFbFf1O
7r4ngJ6DsBL+uRiQAWsKrELJbYoh9eCAgroN830oX9tsNW1tHAdGQBGZx8NbV0OUN7/f1/Z1wXca
IyALKflq8y6aid4n/DwUB09MSxAm9V/3d9/qNOHWs+pVtEHYnHYrOXvvCH65D0tdqnuPwpISyut0
fCUF9ZoE0lcQ2Jbv+3hmevLv/ZCrbN1eOwTMm5JCMd1EYyTW3sxvUPcv4TnHQj3hlZfxVqNeZjU4
s1qMkSYapz/ZsFFNKAS0K9VLO5cyd5uGvNzXYxX4+dKYHxE5bQ6cu2DYhfXcy2UXyIIZVnJ+dJE9
/tFjmobp1qoRMxRp40Re61BYfDh2DE9CEFYJQMw11+I/PGmOiA7tXTnZDPQxN9P08oKpETLxjH2Y
XPkhlDbKlNBixU4NZC+qsoDK/trYAEsHM8nHMBjxzj76AB8nhanZ0ECxUWLPn0QX3vxWN0mmMhNY
pYoUcx8jUJfeEvkyt+K2+QoWRHVfbz7Z3JGXiKmdHV0mzESmAvPsTMjjX+B4axxewTp8zkMRDBA3
SEgIELW/lTMeLFLR0VHyNQw4nJOic9eBcpRwPP0wxXpCis3L0UOi03y/NZIvs+rcK3VpL9gxbMEI
VZomogo+wW/XrhF1ODFifxcoHsZFEXf6xdGS+fX1YMwCblnY0Oyf9eoKpaQ5Cd2/RK8HGCXfTvLP
3L2l2HGG75pfRhU7ALMeu9j6bppuh1qMWoAciAF6XgIDd4bv5iauycHrWZ1YtfoERVcgM+0nRJwW
bpwjRVY4GAT2zAAUJaTHbtUBO3WK/rEoNRMvNcCi9rayZOBmprOi8/aXwDDNvLySHCsSK7mH6n/I
sgZXKToe24Q4HM4vebTvFJy/8h8c0LbvUBQOXw9Nd29/fCWALE2u0QyoGCANDfsI+tT+hGJfPONz
fK/vWybDOoy3fOxR31/wz2i9Tte4S8F2uf9lwFZSKuqcfsR8Ryoiyl0R9JcnDCSn2nktuKySO2Ai
Bh5EKvnug1sC9qqRpEs9KfJdF2MHjiDfUcuWRSY7dC5/4s3Gk05YMNRZqjbgvqCb7urJ7Z9H3+eM
9p1VYiOZxIsGgmxEvTsp5C5lkAX9m2qng2vpVR6Q8SFT63roGIaHtqCORi0XdNheqL4FVoW4o1x5
zwFHOXTCcBtAW7cfUG/HkrWHEKcdj37AJe5EW6iXK8+02X4TpLERtdfQbyIQLtHiOrGilToHr7Ha
OHjwdeOscAc+kQefKIHpZ7++c9TB+BUtOFMUy3a2onB0JkEh5F1zkpMjudMlOEpDPrAXBkSonCmt
Fr8dldrdZR5sKS1yNowRJeRWy30OmdZdxqnyL4mBkYkgwXsB5oH/cfqiF6U0VHRRaAn9/2R+MMpY
GO48pcrffgIPgdVgOebJTvOBy5TJHaoCMADaRnK0QHfD26v3EoEeNdWN99pej+QeGGGSF8VSdhGr
+bfjv8crcaa0+DIfoENZ8r+GyGaBUey/vbMpa+rsivW2omv4B1EUh9hpkBuRG0IURuQs9Mm81f8k
bVCtiXUjUUkjOoNto/27n10MryeWj1z0yygOo3vvnSOxaL3SSv3105tzYB6MBmqDCsTbJs6SFnqJ
Moi7YSrMmy5q2RHBnCjxalL+NwWus0Fo+B0QR6cfZeilhMCjmb6LWlkRriDZG0e2/KviEK4/04WV
y1ytOv9nD5wEz4dzP3M4b+RGQasR1Zl62o8eIg74mubwQTbzhiKeJ2lKJojOBEHTkQTtGFvPvgAI
TNnMAGTAaXnAo8wZ+S/n3vPKpnOTQUM3F30mDGbLEILQArM9YOAWUs+sw0moNoVKfwSYLBoP8axA
m2KylIC9LkX9wl1Wlz55WSnmSO+4ML/XIWcorpIUN+o7cPudfvh/M/Nl/SjmHVElj0F6qhiSCJc9
cHE9qwyOGRSRTJjyzSIuARGR600PtI53IbCRAqd420FBlcbewHzgCA+d7gYzecwaJQ9OkLNxv31J
P2tPsRyzroDfBVDcHquaG8d6FSYEuIjdCjpyvnV3es6t/GxRmlIrNRCUVEPEJNiOtcy8Fu6VKPb3
dL1MyolV7dR5PIC+tqNBk6u+fdk13e62wxurOe24clAI3RlIjItlFxvEDWMZh83maPyDHHSkoyPC
d/uex2nAvERw8oiLwuoj+6gb5YAbKLPMhKLfc/AB42giGV3Nbc2dJq1NVGYPpqze3R6LQJmXsqTB
8VcU5+1Rf1NAbCoRplG4+NUTNtpQhbkZKJRzzoQpYEc2bCWaWOUqIPAI7bbzV0lV61LfDztrxvsG
HYCobvVUPxT15UkegyKeEWqhpTjpx0H8BlHLemI08hcuANyXCbdBu1zcxKvqPvAK3tIGd8bnP2iq
UrIPjwWDHWy1kQxDn15ctDYmCh7Z31l4fvWXjZqnah3bjEoHvpXO85EjvqP1VxAfGyEX8z3QVVn+
diDibgLKO5FwldbOV8a4JU0cr3uML/tfn91VqkWJ3YcBGNyzjI/BU3tbBw6b4F0NqDrqMzyn6kzi
fB24MhJR14icDE2ysjklL7Gsj3y5EdMOA1NyVGwaVavnXuAHAA5G208fp3B1DTaDNTjXR54uwBbk
3elvFmCFefLE6bV1qFAWM8G24X0pig53CnTj/p33xZerzH2GH9INEpPpEwhEyFMK1VCPtH/P7j5h
k2h65tJ2I2Cixbgh+Q6YeqANYrE6pJzK+M3OzsC7Xc3C7HOesqSNezpWGWC3oY/Xq+ZbGiMFCiJ2
VpGFmY9/TYjZv+6DVhN2vNBzaHnsa38WXi4ZsxP19nzveqYIfBIT256BfCe/4hDeSLhx9RcitR0i
MliEo4agJ5yKxxb1RH10d4gKF6r+/a+VSy+fbwlaeugBrPw1WzHyWGhAUgo9asvH4P087c9FrQlR
zI+Gmj3gGpttjl2CIsITNdI1YmQo8xp1335YCcjhl46ZkJMvthmBLPPv2e2qnwWB0C44zTt+DJ9H
RBUkFsEuQlFW5t/eYLCg5CD5Bo70yCY3VvPaS3ivLkQS4ws7vU59OraWGJ/S1FEM7woCXQbJRzD0
Maq/dbXcBJK2wHtnXFt+dBKCGCdaAnVStWpgPpYPp1RbhPsphN0aPFV2XiTMs9+I4fhK9r1n9+zY
Z87idLc9u01AvqL7JKTZeCkwa4HX6pY9ZPI///KoDgE44CKzUmvpOk6cgsCb0bDHgYP6acTU62Pk
+KUefbIT0vmMcRDlhId9zZbeIT4MZ6o0yZMbUYsRKHvvMqSJ8EWROsW3GbqMvl8fruYm+L9ctfnR
1Aw0VOMueIUaDSec7RjRjOh+GOvtPfxjFHzlQEQnwIt4lpfuymMbTdLiZTnI3/vmrzW922SUVO8U
eSpsxsnDz+YIriim1wieni+tiW6zLG40/fzKbCrPJ+W9Saul3TbKNLh79UZ46P6hzIU486beQISI
OgB1ExLcZcYBxC7uVVoMACz8taf/yMNX5NvB3CHJFspRtSg4AyakOk1Bbf2DBRDxbiExgkTNGBKN
djLzHNpju/aR4xqskrrujrAa3oopsmmmx1Z8HOAaEEBz1NXLSEAI9r5e8ah5CXbmGxve9Y9+7E0S
6Af9BmYUi6iGMmas0aPRtVgDQmdXY6h2PkgdF+XFBtg2nK2AYYYAl6bi1btBrxARUNj/OXjDb0Jq
iJoJYzQLUm6WgyYKMqPmo6rnbAYh/HWOUercTeuMrTWwSZh+Jei5cfMHxmD5LqimFRpiG0OFwiux
nqPOOsbhzv5LlyfQH03V2wChC0+J/85DxcwU7LgIRWpRdZfkBLDRNUlWnMpHy4lbmBJl9mCaFfbc
qlDLT/cH51G5esRAW/P9SaGyJ9lUNZTRCBt8Pp5SRWB2Eq4eh6XtRPmps+/IBghuwcT430frKHmP
9MvjyYngjGScqdiU26OWjSQhnqZ5zqOJyKE0qxerHh8FPlUfaey+seoylmXfcJKdwUUiHkkGIjQj
+Ub/kC0YVoiKrvEG2GBv2HqQ3Fy/Funy6jzI+4K4HxpGbuxVDKR6HOeGewPUURWyQXgd58D6NLrU
p4TWEpM+hv2fsDxz0ELZJGVLsLpNkkCeb/V6TvHxYRkwR37Lq/LlEpwyRyXhI6evOpv3sKnv+nXs
wKSET1vyBNvKyX1gcmnHMdHfeTlKkO2E+xanCIGg0IXcraWWL2AtiLTIermogt3NbXMLQ0bfhs/3
u5dTqcSBVaUmD0FqD9TnKzESTpPYVRcosgL8okg5+FvTzUDyYc3RJZ40C1J4c0n2h8Sag62vImcW
oDdpF08j+gM3OszCud88sY60Itf/YR7PuVYXziCkd5pX5esNS8L+l7d0/OK392Ppe0H182se6Sdq
ezRKFEJ01ycH/SZo6hGIWJDQGhi0s6grNoWrhmJVcCU9ZRYHFwoApoAC3ecZjQqLeE6xXu7bBaBL
f/Wmm0dyGZq+TWYdWAB+znHam0LHjO43q0CsfFQzvtBxkPKZxyolzGWWX+H3dmsCqLmCixZ4mu/j
4dazkQ2wPVreANj0S73+ftT0DLHEQaopqiRz42KbPnki4idXRN7Oz2bMQTOfIIQR7Ir3vvo4oRn0
kWVVgv/TCeSiMgg23ejbleJIXD5owuu1JHmR1BLcTCFJeH7MFWMNpKTOS45f6LYIY5d2pYSFNwrH
hE3Z/E+6PDmaWFBTPNxef16zl9fQMUbYrEG/QDj/jDN92smirXRSgpE0YiJL/Fuq8NNvrblZnoY+
TpMdm3hFvSqWI+1fyRWgHAkq0rIwXStY/9139tWLVvWN8FsW4cgVEqP75GohIzE5E+23N9LTaYT+
y1yKgS7Sy6di8lFLKJJmrGibcUBc31S7cA5TDZb4RevbUh7Vg3kqy1GEU08txDnAE/66k3YnPI1z
7oo7wgs6tTs4ZoBpr5XgvIJ02miIgy5M1QNM/TnRLcJ11CjUOB83efPWZCAFhj1ahSlCTsFJFEUX
OqPk2XmuESZjoLFzRU9pPqwTCZuoREUoKBsYNo+g9bOFxL5b0g14ZHZo4NQsbwgf+oa4wvVbX0y6
tRAVWSU9vIVBPHBLMMx9bS2U8DRNJKK/GXok5YHYDennyanlOCPUpIb4wXuzHyjpDFWYA/M3AHDD
BuUUJN317xlsPl52mtlfMZ5AcAkTDDprchUrWbMZIlNnbTeqY6VJhxUWQfwsS5/K5Ua5z9Ra4Tx9
YTJenk3yvZP0oPBBh3xPwxE3lq7Vlt9pUeEiOA8ydBxVmGiNU2f5qhJLVEaOZQcXBdOmJ1RoXDAc
RVwwZVJpHJVl8d1gSPG8EB5wtx8IzNX1Uib9A8ZT48WUzQW/bHuTZK89/XLwCZxMfqorKEihz2wh
vpw58eNU1B5QdjG1J7shlVy81IBJIFUEKsLy30d+sWGj5hwzcdw4pl2oj3cJxVYIJss8G1glZfKd
OHli2SwSTsjmSoGcnIPBCsqnV8qX9VEI2USBRNCS+PWh1GhzAVUWjjUpLdwXNvZeBxndSuVS7aM/
SCPoE5wZ+zu6TMrDaD+gFSRrfR5XrDYk0EZ0p1o39fnMUy8DkKe8KsW/CzJ2/ZRbzcq9RrJW3xRs
rvfNTk2h0aHAHF8Sn6QFOdqNQjkg8gydCkPKJEM4dGt2CSbpaj8XL0bQF8nNlsfGsj9Wi2HZeRmJ
QsVT09WoztcYtuEX2W1pSUUOdWQaDtNiSnmhjs13ODxe1V5x7vbUNlJLbWMP7a1jmG84KGWyZ/yt
ildtRqpQy8m/H/UW4PfoR5yN0Sh961eCXKO12C23m8xFqZ64WlmNAMoiAJBBXVGZzucHgsVhx+UW
OlQOZ6KxsIiKBpb+kbylRF7spVEKlTpdmb1ywu9yzxDFonBABEJZC66bjzcn9+0g/fAgslDdqe5c
hL0d+D8hoSYjVYr2HBq30PV5DJxLRgm60FpYe9rQ5Z2X1UCQ943ScJboAOe+Zd21U7QXOyYP1eAf
Z8BX2IvSJ1s6hiHkXSWHeJso33V2cmjloZZ5sE5V9BhUtB8ZDwmzhPaFG90HBRvKLDpUmw9gkO/N
0PwvkD/y50nTHstCQ2gF/9eezWXX8UB8omXXkvjfXJMly77ctFhhNVX6CsvgTIqedUhQJz4gimOe
tyf6fw4qIn6V9DHCK0PcC+VGFqMQ+NQfcL/UsByVU7IcUig5zb2sDFOx8AX9BS1APTrQRWEjb25G
m4/uPN2hnPTjIU7R4LW5w1myKAqsmz31GedWfYWydp9DFY+byhuYxW2F3Fv3DusaxcHgEgaqCdAV
akjBv6NS30h0m21a62kowgGIdozp14kRU3sOVPgZ5xqpTt5WKDO8VL7nhD9ymH5FP3HkaQ3f4XMH
ZtwsJ6QC2UxB73vJRqWiaPbmR0ee+RmvPP0Gc/iF41cU0azDrliq4BPWOChKKfnaB5SDobRicJYm
ypuXmP4Ja0xE+dvT9j7igeN342VGv9cCGd5GJ/sdab5uDsRQ8CBLNCJsSDGr2ncwtLpSEBU+/JLo
cBpsL4Gbsjf74ypWe2hp/AHq6fMHGgrdiZAORLx0hD8H/+I1v2V7iLUyZzfNkviq4V2pt2wB/GLE
Ds1aQKG2cBaYR65rR351z8lN6hApT8xAv7ZSEGpIa1vFB00m8tt41Muei6bbHcUNouWpvTOaS3fH
FmkXkjSANaxXSa5G4tPFSoVRkxrM5Ivfq0N5QrF8CuLXwAgZ51mrpLeXrk6pE6DJsCyiGNfSbWRh
uqR68nuDpDynC1S+cRI5UxBXXTmRYI8U4EDsW77w+1JUU2jWRSIpcHtETcSel5kte3w/BdFpRnAl
Fc62IoDxHFAgaXxFbDieQL6FhxXCI4L4x9MdyOxAgO+UlBHeJtPw/J5+hlynrxMMm1b1Z5aUXOx+
2HxSf+tSvHmaj/fi+VuIRSE3RgyhaXJ7Yz+K2RZmAq2fua2LokHo8E5tJ7JmIM52fBYogH8EVeA0
HZlay0xU07IX/BJx+xo5DLUOm9iv4pbE7ul9eEuxRnxI9AUVXJqb85s/QoC/Cqte8Ka4i416Hkhi
WrsyTUW83O4krEKrPnJIhkou/Czy84vHm75sv7cuTsvB1AkIvkFK83NzXxJ+RHLMP+qb1kNYC0kp
AUMx2h3pmenN2JTuSTVVXT4Oq3pRD4N58eLzBI+nF9kDIDa6faG8OWE/ZLUPHyboP1yrBUK+ZjAC
CXmkw5fkXn7pEREa9+YHxBRg8HkCGDDuJQyEJchBfE7fVxezk2LlD3tx4EILz7BDqakggJqpDbRt
84UrdkE14TMsRou/xDTmkjlL4lGF9ENHZGxMq9dmbRoGmHMZRwq2gHyu77Son4NqTSjwtt8ViDfQ
epCCRdUIpBd/urBHA9SRmFlQkiiHlvbdWy7O9bpHTC1JHE/f4pjk4U1P9z8CFIf4RebU8jJt+HiL
RLXcf0dqu6GafT1U3aScum0xedAbZWvCdzdoZtD2+863lna5BPUkpXqeVMRg0kY32f4+B2aJuDQD
1huPIV+Q3e8T5HnuMzC2FgcHa/WJnbrv5c9REV62OwpQUtB9vyWZssh1R8WkwVC2FCpKi+OZtfDK
4J7xCqZHxpuhi8pnSxeOg+PBtqrZSY1JSPULQS545L/Cn8IV4LhcyyGpDl5/uREKeuEzSnL9OokC
6DAyN2ehTCFhS7+7S50q9N60WvrWyG+yH9VEUvGFD8kLcgh4U9sbAW4rxfDSXugMF5Jyjo/2hy4x
oHAxgtOXhL3hDj2Dncy5JbqNE6SvnO2Ja0yAyXMa8nxrFaK2/Gur4D3cdHznaq859AhEi/f1lWyy
aubgpT6ULarBTfAeaHa+SQYPUXlUfp772xueFuUrjKg8xhejWpvh3FC16XcZCW7psPRsBeReyqpb
GmNipHYNPZLFo2/COUD2/T2N75Uc7d9ZFgz5iGNiO0L5R95lzUPEUP3fAN6mBdJrnMEwwtY+WQz6
/8fyiZu+Yl27jz1+0v7AKfSBROqhrPjFNEa1CGehuTlkVC/obJT1ktcXz0p117GoyA82bJW8FmP9
6DPZibVBPlsx0kSnvy0CFC5BKPBLNe2RJHJCNUsqmGQnu4iwpFRmp6QD8UHnaaJyKB2aOjwCF34y
wklmQZYJ4Y/s57yqs3QLT4z3xu1X5OpmkWlIYo36C9kILzNKRZDi7RUTQm9nQR8EuPZsLke9mzuq
aexvxP/UOJPWfyvOB3Md6+wUjmNlOaE7iKtLpYCsWQQe2IlL2uzYlhEUcjulzhZLJ3M6RjI125T9
a3jhc3K7yMm1NeKxwCVPkhfwW7qp9cqRwnaXMDBVt+RZMqDM0Y1NvNc+f+/ol6drIcQ9tIEeZEZP
5o5FE6I9TqssDc678ppHMjvAcyr/FOnFHyS4Sh/NmQNScslboTCjXN+fOH1lxDwcRHmpq2TbuIcz
cjAT/CLz3SUbZ1ZWshm6FGeC21Xy+sBa3vixFPbIo2X8tPCAXqxUQqfahWjBGtrXslCxb/loNy3X
ncbxicp9gHKWJvmpLjjFFd29Z4bfubzEx8LrPg0AAfJlkLmOvjm/RVCyaOckHrsw+c66kg89+scj
TSTRtcoMvGTYU4V+xlTJ63n0zigR2keGiXwvDYQBDit5e/EFgctugOG4nM9a1M2+BQtUtR/ISOeI
ca4fxwgD3fs8nQo693kEDubX1/br44SU//UbQfcb+jr3zxhN4Rm9vRvSu612rox1encYPSnR49nD
+JDsGyTIkh2oTX//unbJKOS50gx9/+j8Ot9MKg60F+AnDuRiI2f7GrLXbav9iJRCLkPaWgaxIvhP
dZGBgXuY1hAUx+2qIS5SC4Gl9sOMIEkU3crau/UMy3TelmaDtkT4piq2baE/WxHcopxJpI3gNZYP
2sXi2vK6tcmrek5N9IL9ceiReP1+3xmCB8pWEuuSqRr1ChwOeaxhstb5cqT/eFVdRqlOOPUj76nJ
x1PAJm82UKWLe+VkXRdXZ/aJHLFAtq8ncGWEURldus05xCAZ7xrVnrA/ARoyAt5sY5qKbuLDRcUv
iLxt4ue09wsuU2DRVM887UrIJEoepRPk5L7sGAMJR4B5bIaIKSr+Qc5m7W4HyEKRMw4Qf/1fYyFa
/cdkqla+g8l2kxijJkABbXdV0h8zS9SOjjw8F/NgHk4WFRFiN0kFo88Nj8DKluQC/oHyTo2lDeGU
2JAATltleYUpfPzXiSOiqo6jLX60jND33lOJykwuf3CzViI5euRoTvApeLflkXncct+PcKSb92Ne
JPTF0J0tEWf+S3h6J93PhEia2pk+5D7u7LaXo+WXVltndSne4YMyimkRwBplqqnGSDIyNaNKxHlE
l66FzNd97A+ZeMWpepNaEhKI0w4QtLcKxZ8I4QXaDOiVrPCNetsxtHeeNtQhHAjxiDtrIjnsSlqr
lz31g8wfkxXpDoUyjJmMxrjsE6h+asqimPsu4klK7ebaWEnI2UBodjz8B53CH9Dxq5ttiJiLh4ih
0uaiA1m4fJsht53IVNvjlHfx+1VoqtkHRBZzJ6CuRWR+sK8EEiPLtMT7BmdS+Ose5cwQU5+FTQQU
TAGpb5gSWM+mPDpspRISnNsbcDACOtMlxR3V4115koidSlNqXZIU8sct72PPkYgFcZpmwL/K3Sr7
839XZkYDYKOGYwoPFSK4ByLq6yKuAaqJnm9S1psEcrOYYI6tZ09AXDsijgvcUbqTU9aUoH6Wp21B
pyk5+SpQClYNQ3U2F9IETnfMdXtepOefzDUoVNkzrVHcstB+nK7yuvREIwx74cV4qi2n/wkuxZVo
jH+wSkdjm6+STikapisi3IW+th9IwikJLzuY81Vfs2Og87HGwhG7jT94ePKd3Ixi/BF9ASj2yYqc
Vbs6taw7badcdKsG25x6cc2HB3ojg9+cx+om68bhbcCGEamVwmbqSI2B9jxRecCmLBmPRqFjeGel
++UaOo0jlFS+TMUThV3qSh6j1R6LSTcqs8DUJ9Hx6rOQTlI62MrL7wOS5qZ/T97dNsGZ6JJFXDV0
YPCCi2TzA49nXvPzVFg7gD8VXYPy+DRubGbWTLAx24fOeNP33LH6bOXL2uaQtmzEQC/fa8GwR/rc
BnF9Bdh4A9b/G5lEUUjEzLvKOp9GrT/HpozP9fC2tpt5a74Jkqs0fYWr3itaiJVeFB3wRP4nEemL
QyKxZgSrrY1vsydBnUWBm5ew1vRzqe1iobc1+Da9iptoUDdvKVdwGAMnTdN+x+1/ByQLqQaX4JSb
vqy9Is7C95HSoiSffVP4DZBr04VfnJ8dWfgkw7gTzlLH0uSHk0v9pi8CS1KxB96OXcuPqF8xi9a/
ludTDrpwOlWbiVqUn5xM8EoDQngns85PFx2NjpNZmsc1KU0Xhy3q1iVbkqV1KPsEnNqYNrs22M9x
mWZsNMlHcUtb35TxP5XbslfGkOtuUAZbRvuiorTDSYkbk8DZIOH1U7LgTf+zsaQjnTp0XaKJvLkX
QCJPEnhSQSz1ik4CURITLd0P6Bn9RTABZ2lCdMSu3pJ/UB13UtZBM7b3k7Iq2SbWDgkymr4qHz2N
ESfmuCJDbs9uFJpMICSzEc0F/3i/Uywfsep4s3pddoPGX719dGN9lMJRD6jwmTeOfZBxE3+sC1ot
bwywdFRNnf6t7Q8SHsJzhTAu5sOyyoPUbHDDvlh9txkFY//o/JMaQ0wsrJG0zUT5yE1QfqPHKj7b
kgQpxEZxgs8EIhuiGiNdXo/N2F4noDySU77e+x8hXifxFkXggzV00/Kw5xyYqUZSC2dWj3O6iYfE
fnhFXlhJ8pFwIbx7aFQWL7LFwgYqF3yCSnZdHNRrq0TVJIZpdrUdwt4yvByw3G5haIyEKERro3es
wBj9id3h1D+6ucjmB6yiWmFRedDWk89CyFRMPdOXV7b0/Rr6ZpRF0oeoMzrv1BWH5Wevm4BE/0qp
Edjl+TYAjPgzIDuF19V7JTWvzJymbseTI23DaDLkCsVhDy0pOc4XaMBEcjERc9yUNab7ilTybdkq
gNw3Q2FdBIA2qyPHc9w9ICXxqEj83nwc0JQp2fYGB09GrfZ6Shua/c4OmSXLqpStiEV9N/EVB5V0
iSAumG7uv1BFcfFM5L1ZdMVC8bF/uPz60CoseaiakIHbTYqb20TQZTj3jp0pXjQsMjIUIA+34gOh
PJp+EYp5TJETfjOEyEeZTqFpFI17mdTOUUzxTCXNzaByzExDgqn7+CbUfRjsFlIp34qeZ92/3GGd
9PiwOmqVwMasH9S67AVR6OXjyCAwF00wD15NgC8k/1rNKkCR0QveVSXRRpv5u0+xoVuP4JYvKM7S
3gnWCaLMd66akAhVPpAwqupFTg49JVPFTYp1uYgGLJTTMa1ROEFKAS9Y1wqTTNwRWPnWoNmVk3tL
4Tl8ZiUC0cftr2S4zgFN5BeFNUioJz3g4j78zPG8iFmtmtOgqzU3m1yn5dV1yl72IK6KLLEdAbVZ
qBdPTLFHeu4HsI5Bcv5t6BSX1EvpyOm9OFDzMtb1jP5Rd6mje8CfZw1dDG8xJb/gEMXv7bXUWqSj
jxAMUeYcOPSPipWzvvlmgvwoIEJuyz4iLHbW6XhODXS8Xx7G+HLKRFjw90cj8d0k1ufbbgC1mjgF
85DcZitarzgiEQNWVWXt9Q12kqwIOgBz8mss2eJ51J0JuaA2aa6XprDun96EZ0rY9zNiXDDb3c4N
ArPSYNZGDA7pso2R7QiXT58/Kcsq90lhudHh52lFrlBL/kkCWvxybLvZueXFRS3z7nV1Zzrp2369
XxHkF6acfgfOPQ2MMLJSLGJPEYDUUKaBjhQbuwYk0O7ycqBaOmI2vzsF6ZKdflTQ30IcDv5Gs6Xf
mN1VLtbqzV56G5WNA4xI+iiIj/zijZTZ+dodO7nFAxlTtRv1646KQaWgFWRHShPBb25VWSN0y/8u
D2vjAhA8LqJ9xeVYjk7tg5ryJeL7MH/yq4GXO3T7zIrmddApvi37O1af1xuPV1sZOcsN76019Xok
JSecMZW59LzV0r25pPGCchsI4pOrluPt6SdryT+4Ffaq1ShcoZLNdtdPAU636cOZgtuTCEZ1u69+
yT7sAtjyFTB8c/niSKbHTYPF+B1XwCAbUoh/Ag5/rmKN6e8sKLxj8i21QleQea9ToDEZOR/9Kp6F
sB/XXjllMBLtUF8dzRF54C3wI4ceAd8+FtjCHf5GCSOBrpRvqkMnqrJjxwjI5tR6Ri2ByBBkNera
9rQ/+i0BSXHUA0/lpgQ70y5V7f204TzpzFQr0vytvd0UVvhT6mdrPOGp863Cjyn0T6AYRzRimyQF
Z9xwpBUgBy8dKtD72Ugd2aTvMaZvBvUR1iXoZe97EImHNM7tj5Kau+ZZVt0Ijtq+gSYYGlYYUA4j
YZiROQVFUGeluB4d6USOT2fPyCHoZ4fd0mTm3AHrqYmDh3oOV7pwlV57dFVDNuQzri0RlqhM4Eu8
31y2Bcx+I2Pa4V4rlcW0w7DqSXAfcJJuhWJ9b8QbwnWgfGV1qOll/kPU94H3qD6AIVXMKxowPs2f
mVhuG07s/UK3YMJCf4hV3T54XIgoPvp8LTCpgM5KbSY+Fd3gAgQZPmHCd4SBsjKesu7kwB+Qlsjw
M4JKohk3jQC5oZ1TkJGkYuFD4R1al9gcMAvr8DGcIQ9u6Pkr7RxsPLeNLYG1kJG5plux8w3xM0hg
7UOh6z5ZQUYr99GjeO0u2nU4Ua57iAmj5eHMma04Ob8rewJ3RLNAwg5d1i4PhOcrAvYu417bSda3
KRMfNHPF6QLUMV9VIcOgUmE0uYme7YoJyL2VV2FUB6U1A5vv7JN1qBQsBhTT6gC2oZ0PQSCKgstp
M7UEp3JkTPmrmRLmJCyCfPQTY8Uxf2LvS/eP9q5cpzvzE7o36hdNbnmQqEsgE5uMlr9reVZsCh0B
pAV+rs9KZoy19i4Tm6teDYdcY9Qw/xThJsqdLFq9SwAqETiJ3Cc5dAHNwsNTkDQIeS/NXwlNqKL/
MNK0wzkpFrHtU282WbQJor+LzXsHW9BpHYAoYxohpWrSalScLAOg9BZFB8AMcNIdG9q0Rn5L4jfQ
RyPbCtO3skfsdPzLQDtI7I1oarWfN9vjld7otElJOgO1a09q1Muod/TrCsYOv2M0ddhbWp7vhTw/
9lcRL0MVzV/wqBw5gu7tDvcXMrozxRQxCyuU8bvrOBScVj0/Vm7gCn3EMUYv2HsfYoumyljMacH9
rgEwmlIfQQcF+kztJYSvHMwhTS+53Wbw4Wnvml8HTttuG8i5hx9FyfxfJjsHYLurRRVQknB/38jh
i/JjiKSsniAW8enp5ksZ97CSlhTU5HdeKSGojbbIwsq5mKDvUZNpiy6DK0/M3powZtgD5g0j+jZx
5H4Dr9ptHWBRZzUKdF2CORH65SBCbjfQM5B11pBoPBV+aPNmbHqZpSb9suuahzW5ZF/5NuBUeiDB
88XFZLgfjpdoB6IH1BvdXkBMbXaDg0tRAJrCAzY1FGXOnHZGNcn/skKKDBARARm9hhdAY3qhy3MX
HoxEZyxZNSBm5//jnHX4ezb/aAHP6znqtxx9YwiNxshcolewvecSlbV8XJgMqTzoJQugM/RSrqvm
76rgCtoIzI4t1u2s/phH8vcD8RIj2IcLL26dwP6ko03wlnGBi3U7qxjNxn+iiwZQuipOcLWTWk38
+0hwEirUmG8FgObdAESZirVq/D7p+X7oyirNCw5KRzOe1Hfka8zmr7Q4LJp1yQKcVsGcX8BxO+hc
sY3sXKUvjL9tC592WoWv0zr9sOhJbuLrABAzmq+jrHcWoSomlOVt4hzLUexFC1peGxW9nHax78dM
F1RF5ojICC8rgdhPan0AG8w41YqeeG9kPoXZlVHR6OqG1PlcqBLp58evda9sm2OIbzRmJIUV0NrM
NSAsZFVx9jmJLQhM5YQILymDVD2YctfM/vnKzAXWeFj0sxbMmlC41uuOHcR072VyE9JcIbXseYEj
Hgoa+AnhEOQUzJsMw+x4V1C8S5tNgxaeFhci6QhtoPXRvvi5piNweHlgHZoH+/EzjRBqA+RnKJIZ
0tHILO5buM2SQfwQGO5LoqXyQ74jwjayh/D5cmq20rqLT5A1Y6TXcwlAkBx9tAKBOkvNwDKNBnbg
TtkrYct9amcIhdisD5aAWbi7+Mwr+2HbrqI9ivZJSw05uCerXLJP4nmuoVtRtjf2nXgD4MiKQD+E
tkPWyoEUtVkmRMnaRfiN0vDLqCEiJOXF+577NR8KbIH+NfMPCV7vIVyOcLRG5+pnnCZOzLH52U/+
NcMLq1qK45V25mX/8YKc0433OpXSPe37NBJ5XzZDrFttYu8OU5KXpb5P3LYMH1/LrYXO+lpuLDuJ
BU8U43gSEXxx1biix7IMz0Ok3SkjuZlT5HNx3QzZZ7xIzZ7fToleGTAB4gjteQIOJqd8tRZ0t1ww
yXW50ZzQYJhrU6LR9ytB9o6+DkNvUGs59bsNOo/Zk6clAA+bf9yn/9/r4LKisVtsGJP+R5Yypj/P
T3pdQKQwLu4wAMa83IzgDeWx+BPjU3WWOa0e4UHyHqUCPp3uhM0FXvS59vjBWbKfuSRxIQXhLvDZ
VmvKkFQFbHbCDGkCtLoePDUcb1riKLZMjG2Ak1SBaeBeFsVq66UMIOkpfQuLI5M3o4FXGoWJXhkl
zfdAEaA0d4CkqAjri1QyIAPFO0eT2PaAdK2uq3oSNSUSniNdxGG6wf7K2dcbMzR8Wa+YLTer2won
xFSSSASGwmglcyceqpCemA6KjQA2ZaVx+RhmUz5Ry+zbW2//ELqP078ZLE/UHv2MCsPccdr3spPc
8U41PVFNu8KEydkD57DpELfPHmojSAP4W0xnJUo/116S3QiZaQMDBeb/9LVaGkNYnPxOleKeBskK
Utgpo3UEG9CwOYVaN3QxJFo/np9lciEWtzZqr9iJOOipfOFdneorHxtvZwD9yjbMUa5SM9FlR6v7
Hp/E3k9TRMDpQe69uWqmhLtj5Q3eIve7h/+kQoMFO19GQm/9Pc9TkvJaV1ej2sp8XmHBpbcD6sjv
X/3x3BI/FDmqSeyGnWFhk3HwpOZnJiWRVSbIMW2zHPMCTB+FLFp1bqP0JQeE7emLeAunGrC46BfT
XeiNgwrWVj73+lT8r1UcYWUlceMy2abb4IgsB0MUjrHkFFb1T9y/tqUYuxXyM/bCQUnJqYVz72Gr
AfSNIerEmRcpSyRGN4ohz1wa47BBEW9suzQsQ7a1lWpcd2ZAirBNTmliPb5Dy7xW5eRZ6EhIW//h
QPfEwdydVAdwpNbgNWkE0kL1aUciOYorhQfmPh3SD8QxNxBPYTHmpQivqLa1dQXuc13ZBHun19hs
aFYtda2uvG/PFzhk6TQlmEzWA2fN0o4EtF4PnkmpdOZR+I9y8+UeGVyz0q/qVx42EPYAFTACEwb5
IBPyWJydSCaowD17TH9+a74U/eda93RdX3KmIXhoNVMpVGXMSjCfpPy30iFOt9Ms7wlW3Ap9J0uC
Uo4O/PkXY4I33L2y1lyyxEoCnclzBScwncaRy8oOSk/viYm4eRRnyZdpFdRcuVqB1VHcjnQz+Q6r
WnZYQViY7MNxI9rCuSfFyweiVG6hvRbiiOFxEPQe20UKMluS4vyGilueWNJRmKhEWx42HAJZvQxQ
AbPho1KCaSP1YIl3kGv0kAMh6buPstfprh1saIFxIB/3SvhtI7hBnIGfD913jY0gaihnp42fC7l9
06hRg84zkIYjTo3BCyaqvvotHaMZjQ/0QFiTDIc5/ilAf8cJeIZnDX8BhxOfIWL2FQNM+OZ70/LR
Y6Yga91tqY3flXEdCtOKP8WRLxBGD0DZdJZL1Swv4HJXPYblU3d0euV1AP2OK6H1GgM0jKFdBcUp
1S1/EdCQzfhFxk+e72mc+FYS6XgVYoemXzhW2QVI2omdtOcPD2O6NVlLjA4pRPrdpQdkbxqUU4MX
Zxyx7YgADqh/UCCjRwC3feOHZNC3Ye1bqh+0TCVMbZt4kiTqOKlmaSXauoa3SuKlulHPi2dz3aLk
bWeEWGcp+W3JcPpJKLO1/IWDz1hUItBirIwEFjr+aeAsA+CaDq8RskMVyKLZ7eLjPBXg5H1nULcK
9N09CN0IKzRxt9/hohh5X+WCjXbjGfRhDsFHTAdHo82BQUXl3YlHx/+b1QLq7m+2VNJd5mT6/8hu
vbGS+3AFOx+K8pB9g8Jem119aiQ7LgNgxWc4KmQw4HKJZHG60kM9jjhhr4ik/NasWKvGPRrIFg5+
t7G4NAL4rU2e7D0rQYCoBRzbM9HWIc3g/k//MzR9iPr/lszVXf4JJcjRVNuUc7/uB1VBxrZoGeGq
cRgOH9PP8UFK/nBaKXgSSqsi1iG6wlqikeWpxF9/YOIXtj43h/S43ll/NjmUStFTSF1AsZUkGL3V
L2dtUW2W+OCEd/wWXyKYOdbs6kdYDd6LYMNOgmavzjNHZrUuHbbhWRQWhZ2u4JlOAbjEe7wqtCEK
jP+teHrSIkiB1dVarbmC24TsJHRdxRO13DAVgGC49D4T5E1yK9peayQHHi0c6lXHgV9mSRprTjLk
OpHmz4XVSYm3Tee+xquDr1yjfJEfPDpUQoGPZiUSDfC3JkEhjObhryhukSC+bu2mYwHrVBCuUgLD
fZaKE1DADuB3m9BFZzvJUiVl8jcJr6sjlEIJ4dfy0H9Lo1kgt8wfyrMerpwWnfCdaO9iXWd/M4w2
7SkSp5OGg5L/BZ7yb4F3cV+cW7JIj4gvJ8g80hKu0atlPAvvrQOGX5cVlY1msBcDw7N/l2XVtSeb
RejOg8NJwuR5IYhZZiCh/6nUtjnPKdMKnGewU8ASf8+tPBY3ewNfYNFoOLDHXDoel8x1/6Y7tQTK
d9mU6FTsjcLz9zM4oIll/YU7c7HxtzQ4WbpCcQX5PdBdgjSVsDUQx8LaBu3/j9dR6WSpxMr75We/
XCh2fpuXU6ssYDStVAxlaw20+J4BYgZWrv6W+bWW1+nYhOS6VhCwqP5XIrK8WlsXRhP3eh3J/59w
UafEVHSgVAdVFFrgKxEM4cFVEPNk2NK9UnCUXupSOHQM6/Di0dnAem8yIKNtsG0dyrH3UGQKW3tD
2epz0++lXx/zq6DaMHpohBIJ487amT3W3B7ECgXVtfdqb0Kf+toNyS9UnMURh+/LIqG/W3F4cHv2
yg26IwokFz6mGVSR3ohnxiDooS9MFow99TW7gNZZUVDrYM3KNi+kw1BvDDwYuVaCXPo6nICP1T1I
PPUaF/3qrYzUAgTJAcdQrKQF8NdkzvL9P+h/nsz+RZW5N6YrsnfFnPozSMyS+gfrbIkUIq5kTqfJ
jwUYHaYQWtxpxu43iOFVr/1gXnqsaMfp9qAzgSi6cd/mu5JXBTyYv6rkLGyaIKYNGIAh4JodP5hv
4LtPMiDSDeUY2TQL4wdRTsMlLmvfzthdM1CtUrTvXAV8btrq31y+DCMnktEz4e+hcgGzPx26XV1+
534gA7x3jVDjJEWflLMdEt8xu14eTqwz96qwZcU+8UBDrYfDFXC0XFNnBH9QfjjI0vL9Y4t0Ek1d
XMvYrWqm88DkCNufeTcBbTPMMxO/6EpShZtYBdQO+zK7VAuTCYLx3Am2CljdUmgZN14c33Cwg2Iy
pg7EwzwiuT8RBvz0I21e1idZIRgH/zwsjtRId8yV2wd4QSxiCwMwJEjYTPY6sDY785DNLAn1EBjt
8jlOlQoNblf4RI008PAtn+1hyRGoFVP4AlD/TdOM19K4Yjc+uo4OajEGy31ThPnmTdgDsaVWMTng
E6UElPoby+ftnH730rNXz4Z0OFSMRflkuQa2TCSLM1UlcATXObwI8Mmf7G3vpfSzigT0Ac1rbVNz
8KnpdTJX5FCdNDYCVf6XXM/RouAOvOrTVA0k0h+fYxHHcO6jU1hmk6hocAHMybEv/6pkckZl+qVP
keZIGs/NfxvXTT0Y5mYhoMs9SRpAQ3XMtdXgqZtYEdwe7JqR2mdfBKqoTXAEkljrY7F2JnRAcXW4
LUwWNd6Lvm9bKhl4GdAODuPVmrTcrJhGAP3SnrE5yKM5WCPPaZiTq92UOwoQN4sDKL3WLeRH/a6P
ij6otC1e9s57GhW6wLw8F4pA2yTqwurIbD69R9bPtxNK69z7XAyAQrsH+l2YErNXkYtv47Vh0w1M
WFy2yl09E+n05LowNoqcyuGhZhtV3rj8zDSM1eNADghuDuzgWJy0cgBwwTZyv1E84vJWf+q5YnIG
6qYUeN0cacn1JlQgixyfHU/7g1UjQl4qp5KjWi/0TO4Dm0OlgjAU6CC3yPUhL+9louXnP6r7fFmt
oM7hRR5AJZmEOM0ECsSyDN0sCHnlNX0EUO0P2hS6Z2M1oUpNU4QODLH77TQvugiW64releUtmBUB
7GkxFACnQ+2/5VwAG3ohxZnMiwZH9VsVmLXHRpY/CoEynmp0HeUn6XyHXWJxsi/uxzMReQCDpmht
c4AufoGdHr9Jqrc/rzxyJDM+JU8tyO+9dw8qoFYbS/46NjNodACe5DCrEkUVGHF5y2Nflz4lqRKy
0gVTu0fbAvJRu7t6v6d7Cuew6+FqtzUe7rcE5yZX7iUkJSFMb2YTYQ+QwAoX39s+DwAPu4cSfqGD
btEeAoaoUn5ni8owLGm8Er/GTOYPZc0TskFJUOxgimlTxwdD8vUFHU5KVtXdkoxJSMgY5LD14z7K
XfsZCck8tlrG3ID3pP7WNGXzhEjEqVaXfhYbgfNyPOXUAtzuPhs1s3uz2BOIWvI7HPBuNTczgkPw
O9rVeWbPqlk9MXhMQRR6rEgi9gXsAqqOA6t6NMZSWGLIcLhd+/TRDlBqFshPa7JGX3B3EELiIAsk
Vm+07SjnjFbmaY93Z35Ta4Ckht9Vwr2TnHElIl5R1+XtKRj9C8JyEXLapYl4gFSfe1opbri4dp3i
YcMhH5agIPMe0GqMJpbhPQ6F6W+EBUfKWhoL36DiFoVhYBAmLxbBFX9Vm23tzeV4gXsOXMHfXC8Y
r3eH6ReT4vUcaqWHws36aTio5rJu+IUctiMxncuWgbte866JEZMyrQz2bFlrRqfM19Bqgz2lOES/
dNBTT+kQHShwWhcWAR5AFWQXM3ljTYtfJGvpxkownZrxrbej2RWCv0Vjej7GY0nStMeUPB2OwJ6x
ClPtpZzPHALiiYdrFIWTfAukqdbxk4ACJqCwCHAr1JS38EYQac22xiLno8DSclrsQnuc6MmuZaUm
ZurQQgbhZ5V+5b7hKLK2q4i8lU1e7mMh6v8mLrpUYyYT3AASF3y/xY53jKtzGLVEowxatfHGZtIJ
BXSkKDIT2v9wNy9UUac3tdJW+3ARP/+P2NYXz4hA7AglyyZx5bJklCBXPrKdWc5pYldhWwzDRNAJ
QPor9uRwTQcDq4EQ9Fi/NDelwzlfD69NIc0kRiuGLwxalo7rax+5mBAhZlCtBGI4NMiY259UciP8
k5d1MJ2dK9vI+nqKUAEPSRflnlJscqPsaCk+VZgmELlEmZ2k6LzAG7COGa83dA5V9ekaqaq9pNfB
jTN03ocjx1VPgpPC7acAFhUxpggKcgN1QFttGeCaTscDrddNqz2dqfJ3XhsIcPtOB//OUg+40rmf
mBiwAWKWs1QgC5Y58qzpKfUYWoDZgOid3CoD6d2hhgOsJnBMDIEnmd0hxGqeyepTR5GNcM2BuNyi
q7JQf1yDkBM28+/JreIjFMU+SV+dbA270nUO+SXwegKmF/MwwDVZrk4Nl2fCqLkkXn0jj3ZRm+sD
/y+F6411TpLJj7cXnhy78y0JvklNVfCLAVy+JvUl4t9Xa0LEUkfLBuyctqormjHbw4jqNy45bABp
mrHGMw5FrxWZFBuNwH9xTNE6tdQmaPExM6VdnFS10MiHU9GBLiY26aOR+xdvHWaJuzGrsZhqeo9Z
o8zfJsCHuehISfvH17oZ069JuIp7wNLwPx5LDXEbdeijbIOA73ueXJU58TaILXt9ff4E2CuUtY5r
LG8M8+/9YHeZ0DerFXlprgC+qUFpvELz94UVCoj/IW/cIxMAK/Ag46N6LE3vhD76Gfafg6qbxVjY
2OQdG6gnLx6cE6LCbtd6loSvC3WYny0pmu3KOlEvnezD+b5xybTbZuw+8Z4DtGl/NH2PGRN9GSff
gpzcsq1/cwga+8aQ5l2z/ab9rNdPVd7rzDsqK+ofJ8QsxXHzwKycleevoBSBhozzN0jEN+wnNqBp
NjdmjV/IeqTh9cpFSx1vP+nS7EtiCBcESsRnLui+iJdPgKHuIM9e4VnxUbC9RcSZJnFzxFK5Vi+a
jW7r7SmNGN9Fvmn8x9k4AWCEj9k7APIq0omRlYOgmyH4/CO0WHHurrtM+3ZdSX6m4xN6H5ERMsxr
u0A5hNtIKNjpnF8COZqreDJvivCG/IRc4PE0QgJV8EqaZl0atlAbEI+qYNintZE8WaOctAf1dCjs
3hhSGCa2m+HhOUPDmWtBuocNZDtkIuTlizXu+Zr/zRZ1Nvo6K8CUzCItPVlPiCr/6xf4+neUNGcV
BBErUbwpaOctH01TxPUGmQaTQTfRgBdR609aGU8iRmPdmqGv3klCY8B/ZouqfUZBMl8M3pk6BXYs
i18RbvyokXiicDF8whf9NwRDKJszZYm0a18d2X/H3muLBrDVz0f/LUSnNH4wt8g3NP/7P6RlBEEH
s2ylba1dAr158l22WQZncKwZunLsFT37SquzZMLBa6VPLlOzMOy9HX2Pb8+BX8Vj2OoKBJ7qYSNc
7FHVfdUfRDYC5rOBHMRxsXf1aXoOZrrrNuxkTSpYGMGUOfWrUzgkNHQrQzVKSDfzZ+8wRosdE3G5
QBHkxotdtVgQirWE3HFiWMC4HCIw9mpppxDgvI85eJ2v0H8SwtbzqKUElH68r8WQNCE+hnVIxGZF
d1JQsDL2oFsQkV3YSdUhsnIG12J8VaAQT5VOFAoEb0N6UZyU/is+jpFpiKcpgIzFDEClFn16RYOy
3aaoWCW2ItxZ6UMSGPne2np8dADxcfUY3qVZ7673K2UePKO/uCRVa7NRs/d95Sg6zdu1k7MbtDpS
MsGQYftwhmkTv7bg3TeO/vCgzfnleWi06lk+oXSxoJM3J6cz1AzUChAyHOqyhF3R0MxPmW3EVWHp
YDeTzCC2vl6zvnRmhwqZ2JBHLKj3Y4kWbU+MszRqvqvRHEkgGMZm1cqL7w83SedSzBOMiXbWBUIm
WnUBHucxEUSbDZJpawxpeEAGkvp9eHx4NsqR9cilduTy2ML3wokSAsML+S9A0FZzF41wXLFf9aEn
MwbBynqAJ8wZBKyol/MuqCxAuQZneZFMqfaW6G80fhvLINVYCOIrglJ3siEKcurSDqHYtSD+xaPG
bFcNNy8w8pcxKn8br6kveyzkfwtVCi5h+/ZZmKQBtQMnR7uWe2vConXBKnUqPsnIboGs4kOko64X
3hbr0ClPEilEQDlryHoJs3llUh+g21aUYf3G99E0QuoY4XB+Oyd+AQMy/LnZ7tpy8kA1Z6rKwj0P
i8qz0MJoFAF/h3n9aDvUIt8BVzSFhSbd0bcZz7rxwX5/34BXXdVXX4ZlMlabvhcmp3bnLNMcIibZ
2rwoIIDqIcYew2USmcQis4le7HwKHO1jigV9ypGjvyYf2NpkCCLvy4GFV4KT/pRSPr1dNDSrc8Wq
p8hrn/jwGSzVlYTP48oKfT0Ldu7/dBzbKedWEuuUGc5mNsahA4OSazRl4S3+hiltPgrB+aa9/dxv
7yXT0gk1hXgWlmZ23R9KuivMNlwVcPQKNRQi+a8Bn/JUq+Nuj7C8KbakeLPpEzoTQs8fUENr3fjP
aWJBoMTGupVeBMG8Ku8XzeA4p0I5X6ygEqWK0tdrr80LUmNb2AXlUnWdtc597i7CSNsQSQoYJHMB
nkIVueHztqrsDfPfQPTiTQ51x65UbRw3hXpCAazcTikjGB+ka+BjtmsbBdjczLHZu2skOfRR0hrq
jW9N/s5HA7uvUCeycGHF4VFPwtq6or4tIXzpg5SJgy2tw2AT8A4KCpHkOIkFGcQrtgawI72lI0K8
D/3Q7p+XNVecH1ST8L0RIxXeI+kbh7BD3FSzoWIp0bY26APrURLh0ITzARBAnSlqSnq0trDpU43y
LQRy4uwJ559G/fCOKj+uEEDlK+Ebinf43UUcSL5T82lXI7FvUYzQpnYdooyS/XQJtJWV1RtXzWyJ
tlhxUNncGkKmKuejsk/DvzBqvIA8tqAnD4QeQmtHwmcmq5Jv5Ox7PlCN9dqY1IreVXdp0y4QN75w
9r8aTtuIw34AC4ehH83r9AcrYAWZT6P5EMWD2BMi9U0122pKzCJ1E7wgMrulS/bmWehKogo/CnmM
aRY/FDtA4BN74vbijtivCEbkNPwTGpRqVNqeEMgVJPIzx0/n+E6kqYCBmClPL2RKLI9LoLMXqMFr
ivBlMb1y6rgRQ0yPYgf9VXj9Lt4VeNRanlNRC12T9mQjU3IEe4Q8WusTB0enEgoW7JQY2IJZaJ/a
qVIOxyKMIJDQ0EEyC58UTcdF0vTK8u+dbZeyvLSAKrcsd/K4Vldt8tlDol/xgkm5RUIwI4M+s0CK
J+JKo0En3e64iNeLUd6v9ZgVDXPHmlxsbJBKvvW59IG8bbi+NiAet00tE5CgyTvyhW3rOYgPXlaY
cxNmOi/80+R3W92Lb/MkRr3xvxzNCDUg3Kg1LMsvHk1qgvd8W8guQpUrs8Q08LvGT/30M/dJudO9
RJv7nkxhP2d6F/jwA8BZEkUo48ukFrTg3+iCUpyrJX0YXuGF/IMJg8WVcot/LG9jpsyu3xX6pbfP
1x8qk7t4MYKCrcfy8fO7JZ1mf6IViVkPCkgXhV41Vgfv0+xMfUMirtEPJeOFbEP5XqyT4vI3MEKh
tSr4wKO7etUiYZq7V/9fDIRdPefSc93ABkrSurTdFb+z/U7OElJ4b1/0ApzzvH2dYtGWQDmXD+UP
VRZwHGtRJ13k6Wp98aa8HPMXoWp+oONmREMtN2pmFpyXLuSVCUkKPPxFcrk60cUe/DFJAgW0H2If
TEqF2I3SsHJF5dzI9W+5dYT6YhCz0BGsyOFG12nGzl8wCnqshZgaVw/8ppQmmT2qdzZrO1qPLrwC
G7sB4HYEYnuE/r8U3R1ZXIIK1aegeB0CDvDhrYTbTqlvauuxBuUCjks3z/i0hSNXv2XqbKhnIJNT
NyVacU/OkRkHRI6kP7koQGuHY4qKZJIaq3uWNLSbNpcRsgWs37Lo6a4JWQOHdDKyjzmir1S+3O9Z
P3jmzyQanOw0mQSN3TfuApOlkuvVAHet91MxzuQQcSGW9kDGitFrCnOwk/bmHGYz1y12uk7asQzT
JRFyB6Rrs/mKfnkGqCKYRiqWa9MrV4j0vIQg+G0PypmFAnGPqIaGPydlGPzO2b8ahEHupyV6zMKk
FOwDebCWPJkocMlLPznVRMfLCo5Mv0+9YaDSp4EbM2MMLWa1pkqfGTP4vso3bvnBJZOJfvvcxibo
5hZbMZb/KkJx+jDOgx2yXCEsp2fSWn6tm+/8COUqDK4FfSPHSPxGCVr+hDSIYcF2l/kXWFFis00y
bFF079xv6cGKn0YWUPIMCY5csAG95xDwcxZVBoQ28ScAp9v/LJyB0OIPfykdhLsrcHerD8hDGVtZ
vUll9z1Cugrl5HjgwzW8b9YlmuLxnCCaAql1yz8P0w9bl7oT2OJufHUXQo3GJ7v9OEicVgt4vn4v
MAl9UpjmXWDC6kusg1RKRirSdKRxgl61eEiBNlEBvGRlNip3bymxxm3c6MI60uQN1+5qfoHWUbg/
8c3fiCCdIKS0IbLutq7qEoAdfViznzCx7+R2uQJZnLo0nGukeFLLkbxeorCqpb7BuZiSLMiubgmr
q8+GWC0APtRvhF0SeG6iYCBLdZlhOkFi/acxFVwzg5feDUO1iotI4zmyrClRUkjGESrMJ3vTUGVM
cGkxjYCqlETHmH92fy6tMQMdtpcaxlx/U28xdNBFPOiB7thefpgPYCDKeUOJxc9vbH+++QFzwhYN
GtcKqF6SOTjxO8AxheO33UPeDEKiuscurE6sbkIctGIqHg9axUr1oe2Z/zUrP3U0BqG06tP0mCv/
YW3AxOwOFRH7jhq/NZpCtStG0CKDPnrHlb43nRiR0P8lshr7+YTjN63Q9FLRpGu0MnnFHjc32B0t
aZx3NWhddyLKwHDnlXazY6e9+bs1RPhtG05C9KKRtFhCzVm4BbWgJMzuwm9N1wt5aryBK2MoB5Dt
9ucze0w1VewwA8QVr/cVEnrgJ++M1Ta6+Y/z9fVjjuq1Qc9ZXoBKGc0BBT+18y8Gi44IXP63T80h
1eMo3qyowGscYYUVBa0m42tFD/bQAsc6IQ0J2lzoTEpB5MczdwGOmLJvlyWNXWUjx40m8iL7M4rp
lyNzJJo34b2VdomENXI4UjnAbpNy06ELJ3dtut/XKMgIIhgJ5UjXiKO5lKNvGKblF94JNwV8WpZI
5BnMI4VBPOxU/GZCsNCC9PEduZwsPBiMmLXmDQ12MI/nE2UU9X8N9XoS1ZXSxuVm0eeWov7hlZc5
5DMaDyojY1uHbpBTkyslc8/VY/iXtdk+BEuwT7IkhY41K5K45ZWV7HVd9hePSI1seVR4PRAJQQrw
qWnjH5+AI0TG/L+lCudflwI01rt/AfkJuLccHUWBC6+JuPPwyray5TL6pFZQs1MYJhA8M+t7q7py
bg8mlOTqPRGRTZDKMlIm/Al+kBr/TyUHO8zkj+BROUgDHC38v8WXlvKxjX8VZVHiV2v5wnTlVf8p
QYReSy1Ichm+yzALgMSudGqWGqX1h/18kGDq3L6EO51rG1PScD4hZAtstBYxum+hWWvFlEq2RT2G
ok5FILhx46FaoQDZ8AL/IEqcISRNx/W3r27uWyZs5JmPL0HHflL2BS1y4Hcla7OXnVPOF66NHw87
Q10IHPPmqmu+r+3BX5rtvzunCbdLbWov0Sk9Qtsg+QJOJZ1+6+7htL3Fk7cLQI+7+wwuZdvuLGbk
NkC//a6d0gRvhvj3IQNLlTleCy+H/ZX5fJCYwTPrC8VEl6JMJfNiRZhtRyRQ/YQa2tTRUOQJky2X
B/Cytd766Vd5H5wPTbgOBtidCC1em0cb4cyc7lJE9z9NNa3kefkwz4K/UjDzYEPfsUyWcqfV1nNr
lCbOrEPpBbbICKYJa2Vvzai8+q9o2HtrEEAUQPD4gdPgs+4rrJ2ug36kcR9Z7Tu70n8S6xdR2079
gYJkeAWL3YHwcw3WMabGgU5AnyLg62unb6dZvEwo9HqpeLlXSxQ7vPEK4V9HWqfqdLAhFXzivVDN
l29MSmOmw7p6HBlOh/s42dqOydjwjoqwEEZZ91o6MNKOGbmC0ttMith0djczlgWLOjWuzIPE3OCq
Lwp6W7tbt0QoRtvM3MIIpd4IExPJ3bcuNtRX/NwDi7kQeh8E4uoBz9yLl5YpFM3OHMMYbwnhnz/O
+o2sGaQHxDLa/15k/5zDnHU+qlrMfkCZirbxNlDtS2wpm+2HQ3qpd0clhxpzigOaHcvLN/lP1P+8
/d/pQqdwRIWENdpcencWN32Y/ij6J22RIaxMi/oueuMPaeXmbhHVBmxH3ZZfMkxrIYPlMLNRQDPp
U0hDaLWgCjH+DaMYPdjjZvSlJMdBamJA2oSnvScQO/hnF/55/kMZkdmPBCAiKBkGkIQMUZ5fxjjV
7hSfoalHewANjb9Ms2fgPjOSX5YekE5ZYjO39pL9sIFxdLgPEXn6+Wu9ZcyBNMO8PSqFDLnr0Cg3
+hWEeHd9ljEloK5JlrE5DMxJnNDCC2AodsPpQWXnnsl+RcO5rG8AhdK/+B+Lt5M6gGCpViBXZqdn
jNBaaE9x9UVr2B5w3FU482xtkPmk3DU6SwSYLLpaCjRlvG2owy25kyS7DHBIEL7xVnYJfvR6pVWC
Lcx+k4bBUyQn2UtlCxNChX38dZZQpNr87QukFCHSAFmB9O7bB6wpLVhLvtPniC7iTwd8Sa7aMrcW
ioRzlYFCL2ftqkGKEf5u46ESsfgEGzh2TL9/Krgwju9yyr8ROECl0UDX2VRyniQwEFoTLIXBt7AA
iG2NJUpX/vSwWhOW4wotlQYt9vstoV/ANtkrRZFv9R6UPdyb+3Xqu+vfH/DHWgEEyEssft3M9Oln
Phx0Kjc6ruXhLSyMDID11mwQcNL18gy0wpXEh4SWL3RlSN8ksH0Ohhi1YlSRoDPuD6KWTBLM315Z
0kbbG5xAUe6ekvvxSDPxdhWfF2yJhKuAGp4LD3qrm3NxCTaBoV+T1mQQAYyWfVrI2MATOCFdEYJF
7kwGZus+TlyMyYUB282nIuH/KMgzfzjXUhOcjbKHhukBbfcvjECLZYc0RIf0nZnlTThtNjo+WT33
dQADGogE3eajmJJjz7wGgmB7Tendho0kJZQVFuo8ddTzmMWBQxV0tUmHqyqMBo4UjNM9Hd9NR0io
HsTx8eDwFlMwy1BCiR1KtLW6fWh5sKkftD1G3MtCb/vm5O8bElVmupVQMqTAjyfy2FdQ1pTNEdRM
FzVDvtpE8OQJf+0NgDwpobURadfozA+y0ht3rYPxl1YCG0baSEmR8WzFX1P8Agg2gbbqNqnES0ZN
UjjFBstbzns6GlJpHA4Zg6pm34k7zYQb2sXJOLtDOAD3I483EcSG/IbrYOfUd3DdlQUKrAPikNAW
fG6fm7vPPIJDMHb6suwvW3p3bLLoJ5ah53L8lpZrbh3H1Z4H4Aap545VF8GMS7+CCbqzUfFYcXZD
GzTlI7MsYMxLUwrM0CbkJDC6qV85vv3kEk7MHoF2P7de3U4aiS3AtwfWrrn5bcu8yCKbpTsJszF7
yNxBGuPIw6W8+vupogmpRLwZmVuh6W579nyjbaQZpmw+icfbpM2QlLD8f0R37mLQ/Yfc1oBtnqsl
VhxFabMcJhEcCnxwlvjimEFNSCviBVyRDAILbRSMgS+/vR+BuaHiLbsQska5K8PVGVG6jWzhD6Ct
92TnsQMME7HB6+VTN5nOkJBu1B44ndVF52+6za1MXt+ls6BaaVY8Ratt2cqlWajPsaLI1XS6PNJ8
NO65F0hpGzBfZ9yAnX/eTfy4v2ToyPWFXzOZAovH12CsMc0koSkCQQ1py+X82txfocGoDYkwWPDg
31K8Dgm/vA3iHQSI99BuB2644xzxHyVfWvE7s5Y6gjKUDe70hgXyI3leRUTH559RQueCZZRUGg1z
AYaROr0R+z7C6VbCT3bzWPAyJ6duJj2AeW5WweWUusgwdxIFqYxhTqbe0DCLjigPMEdmB9kbfk/d
p0SmlT8lgUqchjknFRAzwwjT20Gc6HVtNGujg0/nCvKkDml9I+Dg/ejbO8oJ8QTi/RgNgmm/DJRZ
Vm9eLS6hwFt7OiZpGxBQPUvCMcwWwPF1Er00wL+nRb5Tgt9WOdcAZRgneoHxsMN+IxOqIbwzeg7W
OC47Q3BdyYyciEl5zIIEzk761JBB6cfyLupj3G5QZQmvGKdoo+lWOIPdVH70w/Od08mGQgxHSpo9
/8bSf/ZLi1fkOEGIupBDmnEpcIdl518+4rqo6LU58dfcsLI2sxyxEysREmpUVuMAgeBruJTQIhfy
qd3JGiMrsWlLeR1gA8Saw+zcAmTroG/HQ/nErtP2YxMTrtzz65zBywhMjkOEQEij8jNbh1O+RWy/
t+mxdq5Edgt2lVDWuAZZOBimOPbPqa/X+BrP6Yt7mcp0KI3QhHCJHOF7lPQL3XOgfKQmKzYNkwLH
hnqSF+Yq0jxLCtSwp4jQfYO9JtKBChZ5BB7E8V4xhnME7qmZvnqtt0QvfNb39kp55ufcdqXgVjRV
ZV/XNmnyA+nl9tVh7QvWj0FLZgqZ7vassGKGADbXB/unwrDAlmmQFWO0If/vPfUJOUYglNGKYrWN
pP4OQF1+3JGEdLp1+S0TNBfdMefYFtfCgac516qF1FQ9llNh6OCj1IiaW/iBDC6SC6aCTA31L1jK
P4GUHTAdsltK/gPXcbnwEUQd1sfy4Yb3REMD95Ad1Et3kM0sO7mJ2C7NnGmELTs9zJvPAFVMt1z1
SsVS73dNNVDPTxd9xjtO6P3MsVFilbeeiOO8ALmE89dAwwAHV6vwbq5x4LyLlqJ50AI9ebViS8ti
0cSGIVP6p80yL4v9rbqpKL5pXgZE0dgrE1OLs3goZFVzPPpKS4REiPrSxZA7Xm3H40y+tg3/Hzqm
8dDY9QBPB8NQaJ7taabFsFGyXOvXlUnFzE/zkINPw4kyvkEvkEd+KRzzmMi4jBxukfHoz21/xjUi
9UCwW9GSfGpByBuasPvHizD1V28XXuS/B6bQcaLjoWdZRaiL0bcq0e364cBGeFWCitnVL2E4Ew7h
HGIV9OfcxiiyL+3ISRpYIiVF7fgLTMlJ687m5AaX1lvmtL05nMCjF1oITtg7HQ6FwzicuiVPokZK
3Rjko2bqYZ/S8uGFW9xjkhwaCxjKJEWVjrqUCfav805nsh6vmKqb/GSQPcCBUxeWqzOseyhBzqat
8qjbTtrCzh8B5orwOvcRB1UJHIeTNcCAnZbjh6gQGLK5KB9sWHtN989l5TzDWqBA61iAQCV6wcNb
2x8dlLuQcto+YzF7vilMbGBvG3I4Ti977BBuXFqZGzNaQG4d4K06oH2LqunmMG4/fdj1HIGdvgpf
PQWXqBVDEKVXnTBS94xfJuo/7iaFS8PbDIUGK5DqBD6OpfYOoUvAV5e/84iF/llHcj5HQW8mNHsZ
ochDxEYmWRQTeUPfASlIjSBj//N8DxNUsDqMKlufVQ7kyHogZKKzAj4IqWMh5pahZGiSU/U3Z5Iu
kLVWIv5f4lhrZ9+gWJ+fHquZ0sSc1sUWYq+rFZRCTyYMf7cz2c73p4Y9gFxEgmBsgRTATPyuKbgt
QwEId9SDPKjteaBvDGtbqK7qjMPE9uY42VahuIiQs44SJegpWf0qKigdkLl85WuOWErSaPUsz/uf
9dc7lGRQ/M7Xfvah7472R7Nb5/hfbdmffTd2ckBDLz+NkckzSfWnsuA2I1Nx2V1K7FPGglxSx/hQ
ZD8nGlcVuX6/ZEGGARiaIDl1m0/cc+9JFsw/DH1IzPIum5ziowRKF0Xlr+/qFAYmznOI859cHpVb
eU+xYUlUQfoMyLBP/6gXLS9UVzL0lFIRrAIUaFF6+T6IQ0zMhTklkS+UAHsetDtS72MhX9NAMjYP
KKnLIKWWFWaiBRg6cnykUvuTmS5FiuM1yTU+Yj+kqYNAmCU0dPcBSfYwnDpd1z0yQg5fcnApGCO7
6LeyMFksbXhwS5htYb+4IBtW9EjkEblWQa9+CXPK0dC9QGJESPcnJOD1162TVYjUfb5U7r20XjGI
u9pRKxTAw6iT2jRRvBnnWometXqFVk5JWBbOvCG7AahCUuX0j8vCGhY5WDyZo7PVlrmt+A1FTywC
/6intsDUiOPc8DMd/PnShKCzpEKSTdJSpu6dwNwbpWcs+JAESsljqGCVozs7YFkbnmtk3cMTUryr
psLOF0R6qyVCW78O9b/DA81Qgua9XVaJvjoks7GP2mtMc+ym33z+MVw2ZuMJuEiZsXBjD7hiFOoM
7dMitTwvViNt0IrMwfuNYzPWBeUyrN3aJQ7ocT+Q4H9f75mqEpt0Mz0WCF82DSvnTQ1dJKw2To6l
pU7ItIKTI0cNHwU0DvPNdXtCacTbJFHJGMk6HgWI3+5Iqqws/XOF+FGj9uU+nDBPC1rTvi/N9i6C
Bo5wzaRvsecprsq042fsnPGHzkTclKC62M6dVfo7k5Z8bn8U/1RE2T8GTqFb7amRWdYWwnxFWvzz
41N44ynKb3y47t28YgikVnr9zmu9fyfTuQJCO3JY5IHWhr4YqRqsoQerT8ShBWQ2tZ0iq9KBNG7i
lE/HPKW/7tYJ7t6hMZX+a06iE73j5za56A9UE8HWSulJHxA3XrJ6PKzf+d9t0YWZNmN29tzw/DoJ
iUsdxqMPM0PjOsUTfI3v/CPzw3ep30tU0opbD8OzyvDoHklm6Jgq3Dd/0M+Yzn9oGWGIVzgCr3RL
Q5Ke8VjFsLZ8+Vd/HpmvHiZJt3UzImZaeIQzAD8KHIHmPAXYoMe5BAfc/D2nLXkGB6memw8sOOsz
9xZXPM1Ey2slh60GjpHU/0lx/73rRTjMfmezhRtUe7rOlEKrXcqI2jxWCFjERxAJkD05tgtKisMi
DPjd6U5pbzamZ4fKiWbDjeBYjkH0K2BW+wSBlzEk2NO1din3EmehnSTcKERJMLbH7MrHzEpWCv7e
xewaFCav+nDZeihzeUa4CxlFkHbpEWPCvoQIy3h84hbq6c5VM91Am4GL1sYEh6VAFFQc4UvzfkXm
NeiSsWk+bwC+JlcX9EpIjOJiFkHsD2Xs5mrNjs8HaM2gm54vOYPzfjfcXvQCfyzsWBvqjJ3tj3p4
shOlGJ//IBmTsg6R3oyA33b49hz6RclNaxh/YLbZaODOUZ5XefD3h+DMnRjLxNkv8NP1gz6/0gfK
wHLsRHqaXlUf1n1fpFCqKYqJXlPlyCRXDLk9vQDAe2kaTt/mjevhr6QLPulPy12XryQ6AhPDorb9
zjLdN+xSI985E6g+xvP4p3/FFZYbPHMVvNNoJM/UZEY6Bq9LdYV4gGtjhD55StIkEhaJR7EWXR/j
qJ+vHADP9rPPkI+LCCm6qKxPLha2WAxpf3lo6in5jLW9VWh+bCqwy0TuFh8NJ7LxAd9FrDrq9X1d
mffp7AhSpHf97hUwB/MR9v6C+RkrZSffk/UV4ObC+Ww+Mylq1RflvSfkrcOBdUAnz5QO+cPFhg/I
5iu7wj+duS2WLrNGksK/H4wO52rXxjh0/FK3Jp8fR7SfSOktyov2BsW2HEIxZ8ZibhsCN/EQdse1
cY2Eg5Ox1A80Zs/jldK6nv4bMtb0sj/NgB5omC4cPUqQUcX++6ZNJo7bK6j33mJpXLw9khrROFTg
S1mP7onMFr53Y/LQNMLYsJNvvZ8q7iWp+7/oBQSFuRIZRXpV7A935ghTGuHaDLfGkVxpwj1x9P17
JKCGjZlGsDMssC0imy8tjoCT5raS9Q8K9B56wQrRQ0yzOoGGlELKVCYynYE7kBgJPo9UuLIx6R5Y
eXr2XnKgZfQDK/QNLRJqEDYu266mw8sdgAWyuEH3qkM7d1z+L4CEnTzQwi120x8cafn9SK1vmCX5
q1FvonxwbAcZiCxVMeVGDRZryO2j0BACp+jBcwLQNzuaK1sgot6EHjmjLg+DYWTt9IfPS/8XzbcL
2EuEnHMXxZ/XN2Wabwp7aphojTUkY/knBRfd694PKEZcVjW/f6YHEJRbJBdWp0NFYtRfILzFaxX2
8DbbM52L8O5yTOMlBTMdeDh4giZtHi/USXzKUJPY2gQZrs1uXmro1R1RAh3ZVtiDW+bRFV8LUJJa
UKwxm87sfSZhpn4xF7ZuCaY8Wzv9QzlIEjP74WwlQQbaP7E73gAtHeQP4zda9g/oWDVSi7zrfUaF
LeasN+pywICOcAasAA56u0HvlGVnb9rOTAOt8UNlaROx9299D/dGGqEO4qfL11VQX2ocujAHQEH3
qDj23GsNJSxBG1Gb71Y4UzfSr4F+tjyGKpIe57YrPYikDaZ5EUOozqj3aYBZtEwr9VLkyhPyqc7m
xyg6lWfVukFUgmjbGEODQt6WIPqd2yQBax234Hiz+YCsUXGtIkcekxMfFGd8Cec6zHiXqVxUhAmy
qG0isDBT8HyYfWOFmA+t6eU8SEov4K6N9SprmTbN80IeCB2oYFJEp0KJ/BFwoe5PUbYG7FeRFrzI
37B+0tm1JRVD1ZXOcXUfcb1rUt5/QsNZ5ZANfJ4M2ort9H3Gt3uTl7NBLkshCqnnUIBKiWvrVAoB
AcAG4j0Be6Bq+Sl4QPqzG3jVaUg2WNIdb5c9QVgk7iPdKynM9OYK8ThGABRDVU/zuTOK4auGkkaU
pmccaiBD78oApEph/ncZ8MT1cbysJEF7rO6glZp5lsWvhz6bwqTcy2TX9bZNtHxsBfZSC/e9alrM
DN8FXbUnFbCYXe3yzVMiCX0Sf4XwPmkeTY3APO97o1HfiVBULsCZe3ykF08S7bwtO3s1ePVn8ofl
1zqAMsFi/Xio2s96gKR/yRLCqX+FTmpa5wjwGoFJGqJ4n3u6pHYRglDIDXXVIa9XkP1Iaf32lz0n
S/Ke4mjZiwTKtom8aFhhDExbwcdQeXey+/EeXQSgzgZRvmSAkalpDyAF9xRsq//Rqb30Qi2hbxYv
QKKe7/yEFEIgKuIQ5INSeDh3PZ6yQv7M/ijQnY7P9Bum4HfRuh0p0UbdWc9RUrOBWXldRSgDPN6r
kwoCkT7CqJWVDdBN+yuYEUX/MPX/u6CZkw11iFy5u5haglnogBbqKffaF37JHK8NHQk1ntI5cFZp
imJInbObgZpYJuaQ+lBofdh99j/dhve2ddZ5zHz2bBDz8gRyLhLBcG2P1RNPlE5xjwIXSPdzjeWo
d6huWtLBfuh0S5FzntvI2339OXIxcIOyyOjelRIiC/+ibjFKkiO+DWKH/evq44USxA6zFIa+lkpC
+PsIZm5Q73Krb9ArMKRxVpbN13JK6WHGfjVhZhZTXrMzTbzytOIlSqKiU4X0SmPUh26Oow15K5aX
mkllFpw/FV7YhEMxCkVAgKUTdIVXm3aHWg2gwoPzr36APgvDXTyzegTitk+aX5oBoz32rwukO19+
+CBRJJfaafUswp8NBfeg43AdknrsAGw8+FacYmmPHt5I1lHkPi6N1aJ8/tc50WubI44lYSiF5NAT
8rcwHDZtTz4+6Tzr9jqA3HXPKnESkkhSOE7HjhMAYU3zQ82+zMnt9yF2fjcCBrmCPuuW8EkO/tR7
8uy+tsuYSqDrZ+VR6sosHD8XZbJ41twWgxVWWIDJPh0q4XVo5zPnBes/5hSjGH/CEbtgZ1cNWZM1
JPL7mGFgpBN5MrrMXFqziiRugrVEmkSfofMadEjPrP5yHCneYFVdW5cZycak8wQWraKZus/nk6Nb
52R9oDBBtk/M8NluFEK5WGamZHiULiQtUxScPRDmGIjEAxrJkPNGtpJ0VidT3UdOCENHGC2G8Lx8
7i5jrN+ngs1WUWKo+ZxxQwrF/Jq4yGPM6xYo1oLSRM4b6iWQShApu5jZpVMQiqhP/EaCspQtu1Yc
vYEfBrDcxzWy1ZXGEDKWGiKgH07C/oY6q7jPn5K0sT60UIhTrTQYv8P2x20j8yMr5Tg3euy5X+AL
crPor9JaGOzV2h0tJu0/GHVJzbccy+PUwhVcRwfKO0tH7idanU5Lzvd59QjvGsRkc/d4GAXtRf9g
cjTClwiTHNbKlCuQ44tV0HPKlnxeQBmSHKpeqVz7+asT5fbQJRmlYdvNVY6bFJdoZGC4RWkIRrk5
TwPG2ncyi77IoIXZHg5VfDekovkei0/vclcRhmvT6HAGyDBI+foJcpuOL50ztgjLvnUD+9QIXFHC
V7nthHi9rRPjdQSR20aXGx4Qnu54QHA29dMi0wsLYsbQElWLhxW5hLxzx1pjSqPdk5iC8gfeqo3+
wiC6GVEnPB6hWJe3IpfEluOHCsH9VVTQy3e1Xb34hx6z7CaXHKsia2dMV+RwOj9hbXgEtkM88+oT
QW5f93gxLUXA/yBkJkUMT+ZMCbogyWfnjLcMZeuy7FU+MeNZro2TDU54UN0/W1W2Fmmuq2aMp9kS
f/EvhLeXSc2kX1oegeLNifRd9D0nNvm8o6gDl2IsgGw+9KjjllY1TH19olB9DCKan7ndRmCsW3zM
f98hY8cf5p/GfReEY/SXMHb3glWA+m6BGjmjW7XAUCK69AKQVMuxvEViOcWtatiOV4Nmio26HA/T
wrWIItQwVhAFdyWFeax8tLZonYGpbJovq/6wbrj1a89rHr81xihhDWfj2eAnRe5rkaWMdCOXAYGI
gU6FmIqCgdrYlHSdpwFj+A9k4RUq6e7O1uaaoHS32gbl1ixZ0fbCnBUdS4k4l0neQE7x+p0mhaua
tja2VdhH8VI0koXzYB39olekSRP/A5rM4IAifob9uhuZYRAywpV6AC3YF6DEdH0FRS7reZPcBRds
d/2vWVrN9fmdm+bv6kSRKGCygKiTzCSEj8eT12EdeiRGlZ+RdNXJTHw0pb89CWXpkMg0XcG8nMf+
1+N1bKRJItNL1D3pumveooKw/QXbZbLJ/l/3rqfsXdDgZe9zjtq907Schj+WjVtTYDLeb97x+yB6
Vy6RPDZfDmS3+J4p/bI+5bCyLbPkmNHC8xrEGmiPkRA4pJlD1v1DgldeasOuIaeuVVBUdxzWYQIn
mGRmSvRW8xhMenAbvbMOgcqfT5RjckOn3WUJmajXFbTM2A7Pn25hu2BJSicgIBGLKSD7Oe2dHeH/
ENQ65ajwOHNE1alnGBi1vqYP4Ys86EJZfnB7ZHEdyWD5tm2NDvXOVTRnOFmcAjvMqly/PvW4udPV
l8CQv2eGNhu2yyOq3FkdxOMAaOGhnNFPsuIATqwFCaeSjFu+L0aFQWhKUWfMM8JZshjWJIz8kSIu
Gi7QWbmy7u3XUMBxOLCEA3mBYbEGVWAyWeXeGkYa3mpC+wf5vE9HMf1p8XT62ydR+/KMFdPgHvP5
D8+zOkbp2CNHBXXOnhDBwmze2LFbLU1yVq/sxbz5dal4ne5reeJcyaG4hmPeTU0XhMbSlfYhLCpb
LTj+A5EoHuR/pa/hu44F78YJC0dsWGNY0+8sxtcZUE70849bIabnI+fATRNmspQw2nRuqZHSzMWE
/C193ttAV0gOTIzybU1LcoNxgtYFvpJc3PIJOxIWi81BmO0vfA+GmKx4o41Lbkw7ETVcvgZGEbB0
fMhNegwvduvXvZsFZDx1nMIyUlpVG9VfY3zNh5TRpmdeYFmCK8RA4+CT2/yV2iGJgm0XVjuGYF3L
BGeveqGb3CtHp0uYheUoVi9e47Y3cJ6uTf0iPl9L55uzFL2L82oBjYkZZcFzkvleXJGyrcvUXTf2
hC9OCdYBJ1st2iCJennULOieelDpY/zk1yHRGi9ezSctwdPD0ae0qeHs0pKI93HNiyu1KJv2hcxd
QJZbMhosAXyD4YgS6ScaM22E0EX3OiJR4L+4dKJk6qTGhG9qbnN/VJrETaKWfKuuYAEK+ygqWWfi
uah9R68GFCvMLgHLpW2QQRiai4eD0mewcXhgcgHT3o0POOW03OpLGlTgeiTas681l36Pu+bEXPgs
sUEXtOvynvLW8sxVG+wi1cfwyxaMDtEKFsJbWbjwQsIOjSE+t3awNzo/9vZ5n2aRciYzx9YEc9Xn
UVugGOxaFSDi6AiiHDziqaHxn2yNbttXPkyiZcGBXwndraG4g4rov3GoDlKuOecScth0gbZ/sUY0
A55ctomroly4h7jP+H2RhAszR7QEMMzktbZGOfIR1manVwJ0KpYmCTpd+S98ou+jZ5sVRT98DpC6
EDhNGcTnaJtohOH9Zl0IirqEIdYrPptfiEcYsqCkvJ6JunRwu6GhJHZ8nKO6zY00PX9wpBlVevRd
b7NSjgX6BvpM304VXv4msTL+XQ6AZN7Qf9/ZDwhbLir3TIXz3v6w06IZilM2aEksI45qUOyCb83l
wsqvY4z+eeBgmGX26PBQ2tGQZSrMUzAZfOXqPBoJAeOnX7SkQVGR+nLgqYlSsIuXEbmGkBeJMGKI
JZTuVoWq3xFZurtEcllKgV8puf3ekit9SomOdwW84H54QlYE51GFqGE4FS55ViFFXwCchNPoV3ne
LHoykFw98BE5w+AUxhBYltPnm8M5JV47OiahjHF6ptU+pXRPhySjPtvPyI5ITf64x7Udz8dIA7gV
9763K6Abyq6QZ5HyTCoTpR8siEqnXt3B8cFnHaDDKH1CkQNYjn5n9/+PTRWJaefh6tYSFBs37Phi
zP4RjdlHNm1sUuZzL2IxUzIunIF/4f7EijBtgKrZuvfdZVWrDzaefxbwqZjKtsOZUf1i1nrAye6z
DJhJhcwJaMRw7NhnaT4yuOuqhq1W8qADNu4TBKJW4O29+rwoz6lmbKKzsjZEkjotDelCtRKkcG02
4TtDm6OiuVWp6lhYgU6AZ4dMAaILGA7GqqPmGNaw7uc4MaPwMiC1nAnhGx3qi1AhmAqhiv3idXLP
9mFD9THXKB9Kj6ipyxRRnDzr0KWklLgicT2WoqhMTyMMMhqsUBed07+1VjQwdkmtddH4JaZEbTi6
tDhm6GmUX4VBlvFWJheBj8CDaI1VYQzOPUmaZKCw4mHkzgeSGbhBUg6lJP4O+C+LrusqmnM0mdYD
bcTou7aw2yC+Rf7qPdfKWYIfZvL9wrotR0wuIB+4zHZeyHVBn4HuFu9PUzqiFz+tVQnHnZmfydNl
muWcJgJ2+SPGWPQHJ7GwB3/3me/moujBu3VyzUyn+H5o5n87k/89vqzx9vQvbpoyWCvUPHEnVdn7
5oWBKKQUVyANE81+7eS4SrAmD3zjEIG9Z9Q377g7IA166mtwNXmv6ncaeFf3LToqGaEsjpVNBxV6
v71ZVOQLVicFDU0E/NTOJyDjKSVJER8ndHNWKfDFgShogangYi3SeiRGNWk1RzuEjT8b+taYIX2A
ciCGJzhljyy2T+I/h3gTyh9P0udxW6NkU6yeEWOOP0Hbumwt40CW0ALZwix4eKgmJSmOVaB4q5Fn
+M1IM6TQT3LTTuSePPNW6oBHvVKXpdPMVnXS+Xa2FC1J3mi2x+nFZ/VCKL9SEN8E0Qq0GTTQ9xFd
OrUZniSOi7QQ0d1TfBx/CinH9ZZ4TbgfnvARNFFbU6c3YzeNzuVXKhqYp8tF4oACzDPzURzVQtns
1T+wj71CEs0t9WeFWsuIQlle/nGfUsIzD4H4omgBmJjwJHMZ1P3/w7Za6KOIIu9wZ4WeZTtf7vFB
TbfbAt16Ra6xrSNTMdWO16cM2YlNmpyEb2Y3R7VdOa/zDVvoKb+qbYS/OyIp/34YbDZKgFoGPlIR
EOwUwK7RY2qVkHLSEYxFwv40Qy0DRPLbeKuszuX6vDR4DoSvGmikrhDy0G8KcMu3zxbuhDQ4BkRk
n769LQB8GYJ1z97EVAgsNzj60SxQpa7rBSd32YFq89/FLzm9TU84N/mm1Nse8UDMXDCFZsrYRlac
wCn/A2GR0tPcYglX3KnNHsanUOxj9BAnr9ZgN9IqCWG11AlIt+GZZ9G6do0wsK66EJc9ZVq9t8G/
wYmfAFK352ERAKDl295EH6uFwCy3JcpY2oGQPG/HSOtIZMBw7hEHgSzUA6qrQLHVCm9vIwNzClHQ
lnflUyN8abAn6qDRobmt8/NZCaLT/Gw8263KPr5r5k/fndcMO+8wzIuQ5uEH4LyOhmLSwggGQ/Tu
ELZsYOv7rIsuZwri9f4VjIMHBwdNFcCRBhp8cCR3W6/Il6qEfQ98XFolWqTv3d69hszKFxKh9C+h
YSTAJUaAw2vVEqqHLabKsaeCzPhh4gwjS9sPZEVGY81C0LNgGAbn8WASydkpP2HyE/lLkPoxOQCi
MBagXNbhWyj3YSXzKBoCdqIqPiYcON/TaXwgIyw9hDKGRbMBUmhkio4EGubMOtOT8ap4gmlsCnAN
Z7E4YF5RQfyLhc8NyKh4kFurN6VYjB8Y9/brxIIFnDs+DoLneqnswycWyxb1BEq6jo6+kXQ8kKVX
O7TBkBWdfpqaNY2eSoRzuLlyjX+ECeoQSSeQBIMGTWwqfa33xiR//zH8sONo1P7pcoDmdRDLiXZP
k5UuYxfU9PEMu7f2HX+/9KSFR+n0H8U5bLrsKFFnPAUxSNFRW39WQr7fLNYQnGbF86Y685Ah1Ap4
WlhepMpMbpswNasy5fTaW0NsBIkax7x3tyug3DPNM+7pIFaD3fnvghOb65cTe+CfNS9qQL9K1/gK
wr3lgj8OODgaR0BCU97svGqaWRQakYcVi5smbAXY+uUwsSSw4RPGUuEsvs/BDpylegavjJtm029g
dZ9L1jry/m+O1rvfsLZeOXncebOIHO1OYlqkmwoteJMbGr08J+eYfNC4PaCv3R348AMFdBGetPAe
z6I6C2RF7QjM1Dd7czsWYRJhqOa56L7Rubg5Jq1SgORG+1VTej06Gm6eV/mrM7wkFwYKFpsp1n1w
bv0/k076mQaLm91H6U2BdpbxjR/JCEHXAONUI1MVdW2X046U7Heu4UMmBV2QsIEFhW8oCCW8ge4D
yqH9Wx29I45iEBiXLiohbXyqPGCLV5h3KVRT3nKLVFtPCXJkdJc1QUPtT0UQYEqHIc0mqmbzvZ5e
uBl8kz5BQqG4I+Qlv2LxK8IcSwNwb75FNWH6tTI9fXYu7/vwq9VQI80wQSLeUCly1qM1035uwmzF
gJliMakQY0wpdKjSMRsRzDf36mEHnE9wzbOKNmV6//8yRu6EpX45mpPySVNuTD7PaBZDy3e8Kbhc
mzJnxdD7yiqzlZ+Myg977rDsMC70sLT8zTL1tuXWQjOVZWPxg7SxmWQ0V5c1aH+kdbC/dhWaWfM5
qeWjPXoMldWCYs8VUHkndjVEGtmDW3+CqcTVkJXE7jaBEjaJQ2nxjtOZrdkIw6Iq+enyakP6SUQp
s6fMDL0vApFtnjLNiDVC2mTVWzxsihw9ixaMOa/TgHg8nAkH0pLG2wsQ3BrUmHU8K8cCFOZaR+CI
zLrDJOpRUX8DcCCq6ksSuJFBsxW1bVjg+Z9tKh9lhDXRuI+ipj5tCHWrEt2vUdjq1QX7mCB/JwSn
i/TP4bgNjK40tL+yJMyDHI98ySnLUPqzkAhrBV4Jkp5RU8rRRkI1uRjKuGEXL2pkoiA3nANTjHAm
PCcmrcs9aasN4KAN8fvr/Hu8Mna4I44Ul0Ijzf7wWNJoGWDUh586Hqt5Hlj5TRWgqN1c3hZ4/rJw
HL4PD811h/Me4yXMj4rPQoWXc56JCq55ZtlUJhFGynz7BDEBqDpeuIrU6MA4eYasMjaBMchCJJ53
WcnjGTr00Zgk9kQTfnHftaMlGi/uCgkI6fSlAadHtbgA0X4OUcVCUk7UXoQS5BKsPxnpSwLE8xaK
DFJZmC3NwaT3wimdNAihV6u38LIftBK8JDfSUX6oCKbcm8k71Z/h8krSY8axGQzyL9ljokBindqz
m8XgP8oRYx1JSKUFA4b9YcXDW5yfJM26664F5PtwThJvEdfVWJY10XTiPYW7SMY1BllZyaolcQQG
eDAL+lcF2k1MWe7H3nv3wIjnq2/TfvykQvuu2jbTRAhpK8FJVy4fE87jOXtnNyP5JHy3A0XdFm8G
XXyqOLiG/rnk/n3lLQtgGIHCRMAjBHUzSvprlYduD9IkhKpen66YJ5o9mJFwXuf4yMHSceziAl+5
hd5/1zt33Eeb1SZPpPIpSheE3RcLaTzqXnfJM98yGBDkuYu17/wIX2Dy3M0ACZCzPLnUOK2Ak/mu
kKNAaLAo1dqB+rOVGVKQX/GuMrUB9uLlleYf6OyKFnQQrkvtRUja0wcDGGCBFJy0hauhLcrDfn6f
55q80dAB0whPl+vEZpGT79KFYxueP22oRycekDPic50m9amWqPKTZ15fQZBpphPauHFcKZLONZAW
rVbFCqdweFjNsr7mIKSoPC140B2dO63m163L34tbA1WbQPUbDNpnpDtQgePoEi9Veu2YhCcfrE3q
5CLt89AaI/gNJVoT2ajsCtyxzYoWGCiPwkCIn4wiu1RowQsSRnbmsf5/OZO/ly0x3++PJv/DbN6M
lXJ6Qu+XkixmAIEvH00TG3G6wh9o91jKyD4oOXmSTYUzJu+Nh1o/ongk8b+2noYbA9oPoudzY0d+
91l9ePuaIcO0HkzMoprbr+LSvuUhOwmMY1AQg5GdNVVjGbnEZmsdP+HgiOXk4FeCZy6GcEwMUxmQ
xjs4/jLWMi4vw90V7kmlbXSyhCZ6DCTW8k5tTCMwX91yaKcQ8BEB7+CpJBa8ogZyr8EvDEfCyJ0k
fBm/gVrQ+mQ+AW4VdBvbUg+B23yESpxiF27rWze/92s5IVV6h9srmqvhKlq7ackj0URgbG6m51vh
6Jh6hjqKEbu/RIx8T1JeG/tme0BEod48ugdL+o499HrIeRNQhGcBsdex5pRPOjeKsV5uncxohT8y
vrpcFnJU7n/4RvpSHEbZ0KevahvKS4T0bpGm6FEHWnFe6JBaWjqVxU5YvjIOC8EXtJ8mV3XLptHZ
sPrjEynpaWrgajWehdb3+cDzSViDYrAY9DkEs583dtIGfcw2dALl5n9z8KIwEswa+4fIF+UVoEHf
C2AG0NdUTrIu80gq0tOnFOuyDP7QEMKv/zDsq7GALoVrMrYat98kRHT9Ff2P1EzQfMluowZLqnUa
AFaZO4C8YTTPM43ldZGq7UDWw3BQr7iHQDDudfbVpg5t0V4Qvda0UHoMRDC73RzUU4pXH+qieswd
QW3Hi446YKwddDebC/rTsnoTjYp7B5ZAXTB+MNF3FwmafUF09W6FYgcaQYKz9WtKuwKfRiIpks/r
jivNYRFKtIJ/frQArL27Si3MKqhZJZJVzbIU9d5yppaBzGe25+Hp903zqvm9R4qADaBJmohlwyj0
/ecIbJpoCIbeptUkVtVyJ5XUO5Av408OeTEjaQYHE1S1ZVlfnONeAvxQorPcx1Hyrxw2CXd/c4Ep
bNsB0iVZ7jdAdKYe2Gul+7RPNgXJ6yWfLpqtO/YU3vCeaTWaEr/GJ0BWTFor2nfMGb6D+7xi2tsT
kd7bS/We8TZBxPtlupOKgYHpEvl6tUd1ZmPEzTgR+H2F0HQhR0uZ3UbazoLiugTYeUxRVbaTOrgR
VRBwPJjIe94SifHF636tJecqQp1mmUQ13mmmb8Sarv/L1sbTMaXecnZr3GPf1yqOkm5vFsMujxSi
bibW4ussEKTc3ehY5k8nJSTbKTcxiqNl5sA+w0XaWlgkiWgGaGjwDP6Tmd8gpoRXJBHBCt9gauEH
qICVMWVsVfkaajyPLmK4kB4XKJQj+ImPC7NxPHkEroxmdYypYJmIhzoDoVJoxnKYjcu/NI4VCyry
CobAT9EVm3lVFQDg4B3BMqTFZWPciQmHNnLqWw345PGkpiyNw1j9YEp9OJ2ziWUioeq5IqciNM88
Qc1uNvliIO+kNprnUGoqMmwY3OF56HM0mC+Ew/hNveMAvpNj7K6kFn7WiwFedjn2nWFUldlNED/m
8in8g4NSdojzyjVaNNCubyjcpQWAycQJfOHBJ4x5VU3PlPVD3QraVZo54yhik9ilNQ2cCvh0N/qh
DUy2cMg8cMYipM1pwldXe5lplJuSWgkXU6a0+I/f74dYoGLQf3l07VcOXQlTfct9r6tcwxnFlJut
hjzajQO7dZWV7NbljDkbP0DUGTzrZT28gZOVZTshjVZUUVn954EfJkFxvAaPiQtEJHCpDW+FI3W9
a7pLbOdtM24TArK2TkVS4lFVhxQofUsuupswqsawsfoP1t36i8nsF+AAwU2/PQrj7ia6F6j5fCI/
LErzYXlbaIXv65CED5y+9GCj5oWXjqhzUZo8cgolW3CezZiDUJv6IisbTfnk372lu87Y6vjJ9BIY
kq7E0wqmz6DOo+NlPj1saYO/ABIGzbbrVf1SJyR7mgvWLM2HUE1CSOAKWqUp57QAkyIydwrxJPJC
O4AIV4q1Yopxn5f9O4yzGSFq4GICdTcfQJHbfNYX8uff0kV7ANKEEYNrnOryuGfyRz5xW71WF5wU
GFkQCPddxd5J/SU6uY7VQJfin4xhdbsgrWkUGLFXYFHgLNolcLgPQWDrNWeyhEE9ECfpa7zPee06
mJQuUKhORwsuLzudO08FhpC+JAb7cbzDeW8aTh71W708OT49BKn7Vhv6bzMQuqU7/M5/BKenqJzn
Rhsut7qWKDDwLM8Gu2gA2Y5WkMxo9XsEycZ9MZyHvBwGmcYyCnlTjc6hfeOK91kqu8KpnccqaQUE
CPdtJkqSwVBNjcmxOXWjjRzzXt1wtH8qcd5OtvnEAvTF02/eLKUkln/awY2Ti1GOXF3nxagynCuP
1D/d1Hcr4qwoydl52n/jd3u3oT+FWyFEgAWTfddZLBUGEmKarX7CbE7E8C6In1I9vY8/j8ocs5u6
87XNlaYkPWsLdcZha0FH50/+9SJu5kngpFF1Nv68nOifb+ZDFlK3KTsZV+6zN/hXSqdOlTI21XSd
6iyoPQGuwq449toj4To1jn7qfi0w5/G35O474UePjEj3AuRmM57TZ/UyRE4pOGEsiQw2N3gFlHz/
4eOYkXAVvPhTpH3g92cnChox0WnQOFR4tyu4CbTZYXy38JJeNKddfef28OAKZvgaAqEZpvM8kYNu
YYlbPuggHwVgsTTwZhgfQ6yunthFQbcT4yIVBMkfhIcm2IGzFHw0QSzsN1cEb1elRpEq9WllLAj1
nEqGE0vDWSLhelhcx8JFNpGJmXLeLJaVjeUrjgtfcO0pmz8t5whJQU4YJOgSQ/WorhEL7LkIjW2z
2BFhYzIgYBlCsIldfA/vb37duhst3/6v8akUhs4Z28zcP9JwhSIa/MoVkOmSLkn29yitWODK7Ixh
zhESTBzxJk/dKFHhZG3JalABZ7nwk6KQLYp22jjwVTRPfJpMOB3Q93Do91Y2qQcTbrK1PJE4QOg3
1B96bK+lx/rxJzduDw6e3bojNAE56FjvaaF5s35ZP9WHI7MLApyg2A+KSWaNZSkCr+mCEQm2Fmqc
BegUYV/m8d8YVO6+E7w+0L3YNrHSWvH7pEBCWBejwdnxGFnBkDCyjC40/w2BePZO4V+XSmfu8T1a
XEPKweMF6GB0k2/y5VAPY+ClgWagkxeL3cCk3PPJKe28o68eEx2Fl0LjVI7ZjSouj8NNHeIciLzi
+GJZsT2fstk8nw9rrM5SGBp1YSQEg60FbKCi+oWb3nLNf36lI2BFnAhTXkrXQIPmhRN92T4Cc5TT
/F1Ww3H/5OOfjy5b/DwSCsgdsNaenNlzzDrX1DK130w+DfZkZWxU2kfqhgurOk1W4ybKyhkC1VVV
vM/auuZ/MEN7Z4eQjE8AfjYiVtwh8DYlS/C7hEAMApe6NRcKhuBRBCF8x/GP8X+VxGvyYp1JKX8K
F/CIq+Lh9JFn0jJJVMbvzq3R39q3uOfnH5XREhehIauLVh5zL0u+M7leGJoyTH0K+i/h4fW1FTqG
AepXFxuZQQVzpXUbMi2z3r1wnasboxr+gl5rIlgxqb04xkbzthVUwfTeOHd+qWhIHwjr8+sS5u+A
I6qnYlJQMKeDenO9THJsYPs+X7GFHX8gZAEYiVrKWKSJNvnofKzXbP1UVsdE+/+C6XK4Lt95lD6j
3LuAxYFpCRztmnIiBar1QPPVzRM/WVziW5FAlEeKdBahHwU0RMKrqBlpytgzOxwYZ6BHjefsD9uI
3IkufAH1aWzxWAmkCtK3KrmPPyj54ik7wD9UHzb0OY1rzNwPsTIfaO4HfutqTiNNDJgLg2EVDW45
Dg7jZz0Hz7qbGWft/HhH6oZDM/HGqd540OUQvDeXRaDdjfbruus3JN4yAiW/nM3viI+kIHKI8NEi
HxRbaYGKM0XoYMnosQk44x8l/E0oZvmG6Qb5lworsA0FhsowgSTNJiFgkdNk8g4+IURdwuwLD6Zl
tyCN0s6y4CysQbclXPF2sFqJQ3VnO/nVAv9bEp0FHYd/OsUzi7VDqYrgVhomipQvrHjshlsBNziO
jItdi9nkwzKH5ZzR4o8x7WXuHVQSBzEMhKAu9mOy0tS9fdZopl5i4IzjsIBhpWBs+owQwu6hztER
JLf+vWGWE/dild2+E06cQiigfaW740aWnWpJbuyJL/FWU6Rvjky/9optQ25NiYqxxGs+Bhle3yL8
n15O3EASNDX1Y3uRHc+hiKRTI3Yszklr1IjulThpqSaJEyuPCn8uUAm+o/5b+hhMQ5jlKzM2s/4p
0+KvRTvqfFn6l0hq9dCuJVJ+0y6y81NmhAgQcInX+tGKQ2WQB6PW6Z3lg7O2pMlJfgbvnji/sK3s
r/FxABHfs8V4nDPkJ6E9SYCgJfJV811K8D0XKnqK2vV62ef/LxV+eSCeatF/e+FAYEwWdBBRgLOl
rcjvcWGpIYXV648Mfk26ma/wDERn0mUQ3ZBrXv/1t38KaK33SGCA7qV4tQ8IaoQpBgmLBX1mc2Nn
oPqUj3hpkrWvQWHviRsHDcon2TVCwzAkZncMsboYoINJaUm82tdzu3Pb/nv5wR5shr8yaeEfVtsr
Ko4WbmiRr3lCXxMzh9P9d5ht6i4exRCIycLBxnx/3OR0jyQTCvZiv+tHk2rtnY0rSzu7nMFXvIJb
CuLKqL0yanNk6UvOLddrTPMrKPJlVXpjYWTXouKTlsBdmFXNq6LT3wrGmIaOE710z7oKRltYz6JM
eGwdItWNPvBNSh6BqwB2vfNF7UXcwzty9Dka76JknXUwj0w80cLieTGoYAdNa8QRialD97pD7AQh
9GOcxD5weG5VJhowLn8XzXh+tRIHngae3VittJWremohIkSsVyk/nKgVJz6Lz9rHGAEj37ZElB7s
h72v4qdWd0KSjq43ZhRksxsHiR0/yObeSq/cevOnM/V+LomFFJnFTE50eBlyOJqKgL/kerIfxBoP
ne4pz7GdHMNrFg36BKSpk/bi1/qI1td15EvJuvq0ORk+ZJ5iCOiInQ4+U5ppfM1G0PwrcOxhn0lT
DizfWQbxgzINwoYZv6gIOEZxDEgfU3Hyp0gIgn6eRxYE4UWltvYkUPlaha1jyFn5lO5Ngx61kets
CpfXmwiddYrQRYw/Hor8OFkK4EzgZ0OGOiiw+TdQyt60+/u/JQ+QrZABNcj4A+gsVkgao8d4CG0h
Y4c/J+gOqwVUaDXpP2bQMO5K4zJcqg2/aXq2vM8jreawoUY8n1UkcALVGWZaw+8bWVKoFHo5nuDz
hJjeQAsBzgXA4qzlHeUCh/tn2+khFub+rKM/jC/y0y0UQzE5J+UdqY48lMknUkgDHVACYYEFOGmi
WBMllX6XmtaQ1SlMRirqWWb9U5jc3EytfqA4ho57As3zYkEyiNMxTHq6Jt5ihsO2hwl5H+xuu5Md
5KZU932QnahimLbPHu+FNUgrFM9Uy3A9XaYgvqD1nz5wCqp7CLXT5J/VTtMc4wFb0sAaA7uz6uOK
PxUHXRn+nPoW2+bD0Q+ojlXwILcLHw4Qu76moA8K72AS6SXDIncZvNn2hjiaMSc6+oW179/xzUXp
gm8F3fMuI7U5zhO8YHxv4ELCPV6VaBO2CDccJPxPsdLDL3kfJwYYpZCj72aGdHZWT9fBCX8dWn3S
NZK7RHFX8BK2EerKIxXACDApE4v5qBY5yOEufHjtg77z4SmRKQvA8r/F1pzURkX0k1svYrz8cREe
CxCXUEHi18RobQ4fCL8RB2Y0/yz1A5loiAdxDh7io6kSA2H48oEecBs8wU0oSOASBDeuiSlGY4wa
l1J7q/sLjXEe71aSWUzPoSmw5vbpIioVzzfzxgNGBO/LMHPrsUAQoZWv2HFFDLOE2ctorNlTYFr0
nTS1DfCjixOnxexRT5vbf7hJU/A/nsoEXZj04JRzFhzUzl4D0sI0i15HFRV+notKmAQLqIBB03K8
C7Oh48l5O/3X+G7LmtIyLuO38sBLPQTCnSwBqgjiKMtHdrW+9Nkq/UQRSOirfIxXqCkXoyExW2KM
ZJ1WL3qkny/gTNUzwaSmwLgOvWuAx+f84nAc7oHx/1zJGb+Pg2LfK7thH7Bw7vqbXy3Rx2MCStFt
mQquCQ36n4jPGvQAqXyLrg+VFcSUIlfVxkPT84TM1UpvcsD7+94CD4IZpAv9NG9QBijc/Frc6nAB
HGiem9jgBFzQ/knFMjq6YThnA9zkzbQi4eRIObdIc8LtAhLo1KcgwxLVYytrUY+dl5kep7uJaXz+
6KtYzS7tNAoV8p+4Y5UXY341BDcAKIDnDmXAbk1Rd5uUpj3B0/qi+3tQudq/B+9P6umGUHTTiX9T
RtbAy79F4zLQRr22y6TyRDYp3U+4QNWVKzqo+ppwHS+RAwJu9cELKaY35wmjjIAjojCKYokxt6SB
fHRDOBbRMcKcAd5vszAx+Do8H7MOsokoVs2qfSkykdRi+qmtajc097IlsvSAwzmh+BIV2nKj0qtj
eWZAa8qN7+6nRY3WtiEqEGiLx3SSy0du102jn8yroFGVUFTEx7hlbBdSI9I2d7AMZf4F+rlJmaCH
o4sKbp3/8T2vYhsuFmtNjSXEBlSDR96KezX9TdqYeQU36U1Ae/ENdRmRpeajZsygDq/oDXbMPkHG
ffKm3OFJndJvberdFMSnvslZQonkbua1y/Vyd+zY1LnvKW3Bsvh2ZCJ79PEaakcnea1R7YwmP46d
ty9AiWdoArbeCQ+ZNv891P+9ploprOab+ytMVSJUWrNdv4iWYc9NsVC09katnDL/qbq1MYiwfkmH
04WAL4eGzzBrNJDVmGbD16wQ+JiSIgYSNVRLMJQ8Atj2nRuqcMTSoZT/7AXk26MofXdz00qk6uv6
zalsqQ2kIylNzYw2AJEFALRxW3US8Hv1DqXnC0Jf4OHOKiKMIWQvCnlOKPWNOUXb2cZXeGZ3NvlD
6SOxA5AOMmniOPjAd3yBgfec5nyI58YN0vUg89XkPgvvVLIA2DxxHbufsp/sz0WHhLIRZAjDvIB4
LV2H+qf9or73btIXhDJkvSzQ51tHG4BWCPERt21014467Y8fUt81eD/lBUezuY0mAFjPyLavxAgv
p8DNt42RkVNkEDFcObh1W9+EFfJPeKxIkgbXNPVGqsbXVfI46fVzSpIDS8P1BA5zXYiM6XrqoyM6
E9yqexSITu9DW50qdi/VJA88YP1uW4yvB8mKfrEpk84fJCtkiIYN/2RBZ0KFOJCTlsOTXH6kE+Lc
sTELIacllrTZwAmEp7nE0Wm4yOVnoQ3cDFId0EyDfc1HG3Mgo2Cxrh0ocNk2SQwX6GXA1G9dz+T5
ewvzysTcL0EFXtod+DdHX4Kxb3rVt97CU2eAddYPFFZIKrNBZOKCTrSQHAX2TFlv5icO2C+AauUH
jaCaSlrsWKOQcf4swlO1JFhCmzWiNroHRPJzOJGP1StpiOSJzDMb6s5T1dZiqLXUkrp9svyotNo2
sJIEff1uJSX2aQBxfyYyuaGNeelhCEqQ/TUyClqMMl30y6hhifNUJNO00ugJRhuBqBH/bf+5oCnw
pys9noGCVqHu3sE+vaaOsqVCJzR5ukuNpwS2/FlZ2L8qDJnu9XwK8FlCq9/SkQUkQC310NhvDU1U
TPEWqvPsjc8WhA9Z+9YokGWYYAUhjgqjDL3LsJY9wWtGGaySf3SO24gRaVpnokzHc1CSZQpBmDPC
gtC56krERLF8yQPNQkrWwiFnQxH1AN7kAuxMEKYYbMT0kylwz4XMuyRlrxxrX38KvF2L073vHJi4
HGZHDahyalNGhtdC8EdkZI0XL+oz+oWLn811WGMSWhfvCBR+U0t3KsJRQY2DvqBwb6ToC9Da4QNi
C/z1NKWcDxAST9Yxxa7OBYP8QfX8jYor6FbDKSbOH5QlL6ZfKIySfBU7xaF48pYzXQleGmeLbhTk
JkFyx4EUWzo8KcH/tQyWQymvQE3xED57edUdcpCbnI45cgaL+lLCbI8Vl8zdZU6AGdfCsd3dQo/M
3QqCKKHgwB/AxM0P2ddXt71OaT2zTlSEzTs70MjxCyFbFXV8DApH+AlrCR6uOie5W3NH5hT1w5yR
UCU70xhaXBE/v57GieD8m/6pAf7alLt6IsPSJgDnbOFtQb7Pr695Q0K5EDqTgOTLxM34k5sLSy5x
TnG+QjQQdhBL4dt5/yw1c91++EGOoqRfO1MDIVCJp7M59l69zN6M2SZnynwg4iVYPBuqAXWKuwLC
CIrhasASJeSWLCVysWUCgUc80hNKYm1uinhFw/rWNCnhAfy8mZkNVjIddUd4EV+iRBZ7QS96T/Gr
a21sGG0H+BMAKdYEejOOqDpwn+9cnl46DOx65WuZpFeqEFcEgtDBqulL4LBlEJKnJyvEeXKDMgwk
zKlFiyp122CtLl5wqkVW5DZ6NnGfJOwjls8p8gxYsk6h87tO4gzf6LlenQY+WrWYEFvkShRkZPr5
1gaQgQ39MsMdXzCZzCFq2r4wAAVtGAWPcxYWvN7TrnVX6Ila5//ZwurEbxHVM6EUIYBjPIVu5yKX
gDEQ/n7Q4BbTlCVOwIKlFKOUcys7Q4eMW/Vl6eaVXvqsh1P4g9xGQfUAxS0DFZVi0viweCX/Jhrc
g5sURerPX/e5D9bqRlmJuH4AzxfEUYeU/yVb5+fKlFzxdFnmZnnTzIdDAtkBhJlHNVzwj1ZwGf/L
+j5nmiozHjfmgWI76+hTy58PWumpCQqOQ4QhjTa5FW2MESooorvHpOEKL40oVilR2Hu35YnrcnQL
Hb/GWyfmre0fLQ0gY9ni9CyjiVca2fD7T0r58V5assFSLAADCtMx7gYMOpUxhzahfRoR3F37quIn
xbvDfPqS3q4AEm4rW/G7uvls+umV/lJ5ajQn/oExpYhIeHx3p6+QucInvOpymJAdDyCajMnMHrnN
96l68Ipcatk0lYT0QLjxYidXNZVDJGdf6YsrKLH9P2XiLVj1km4mSwq/W6bDj76UmVo0ccHbzTSE
VwELYHzZGa4vX3cueIdbhirXKE27lKqD4Cr353apAIIrRkF8nkcQLEwJqpBXNwXp8a2k/eVfjJA4
GgB3JZ/imzdvF8Gf2IQFM6X7JDSlzpoWGhtvf89fLaU2c6bv6vLQlmipmCiBuRmCIa7T3aihAoz8
YAL/7iN6fcQqjVm69jSu6uYSrrSQDMkqV3VBuC7X4clDf1R2oUjEmtp3CfKJEFsM9kIkLYBt/9Yd
2/dpFSWJOim96KU8SHCH0i8qc14NTFOsAWTpCDD5kmAfkukoRI/x0xhJcMdUc9zammRsOrLhgU4m
3s0p+yrmmgxxpM9wgMxmAPFjZK+qT+tJhxPX/54BMWxLJiyEUOMyw/3OzP3ZbvQKAlMuFqjVCUqN
Q7FGQ0arx0dsZt12T4OtxcmF6JTSPUvoMua4U2wPLC3dy4UeSz5aiprGXWwQFz/2VMZQcq1adUS7
C+LqZRRyHwKJMWcFeuqMPx0TBvu2+N2qgbQiQF7djKcaoKitecXyZ/5TrhVOnF9hGQ3Z38Oh9kz+
ErevLV/wvKv0jeXFjwRlTbjxZYTCvkoNqc45vZ1lvFQyQNm9Z1p59BFEWyar2GuWwImZSfFfVXRZ
cVO9OzDRpKLJPWOCHw5ai841obAgSCtcECqOlBRobEWh3h2WpsnekMbyXLwg0LfcZ8R3HbTflr28
oiWdl5BfgtkuVgn417qtlufIKnhVdqlMqJ/4maO9CFShMeO/AOp0PxDos8ixL9OqNMWQL4jXveNz
UM7a6s5b5/XckOyTOrhMC5IhU4Zj3TJ+ahfr7i7KPXMj3y8j3EYmlL0jO1Axn0zhBEr8+mYHnlLw
YhJmfUPcJGGBgs4GbobxVAdXvsRwWFzDDAKVnUp8lHbsjm1jN20qJ0GAOPCc9a7Fq379xUo2zD2A
jWNq4IKUotGZOcF7gFTDjYhKEUK+xi0O+9tft0t6EXqM2M/HLrJ+ygNzkMjWTn7rYUZIwzVpN5xQ
NMuU2s0PUioDIOU/8rfJ2SWQ5vsuIFEbcdVOROt395W8hARbBg12vH2akLxn1cYIBk0hNV89FJhB
hjFxjFHKE9cwSfUyvHzaBOn93kq/438ABTYnVx5HlorfTfpwGAqY9YBdccxk4jsLdIueA4xvbfm5
jqAaFuKjQzxCXQN01sTkcIusDC9FPjrMtUOtIei8iMvC9ddMscMvqcae+KTOS5rWPg+aeYXGTxMU
oalmX6+OtKTQL59C5ZFWEsLifzmRHOmcgbChC1GAqT+/R4a7UyWI7Sv+CHA5WAk/DDRF/mMwNhic
eQBdTgkomkL0phItZZajwkQ70cPvxozloyfeuus75BrqZIjtbZe4C2kQesahkZzVYDlM27k2IpsC
XRe8Dt1pB0DM0GkaHqYUyQQpwvYKNeFCVyp/JUNtDtU0Eoxae7qP+rUc4snkrlvurr7BNePyj7eQ
a1iTh26MECXVzvOWpkgdxnLVP0zq3OvOVqtnptOk6HAx6BaEC8lTVRtQz2xBkPbqSGOxyUBUKMED
0vbqj2t3EYJv49EzNjabh7cr+I/2Sawx0Xw4v0J7LfU6kCh+5b1fiKlDNB3SMAXefSNklk+QFEkG
CdW0QAHySM85sgmfffotlabDXGE92PqcxaRznd+U4p2XpRKV5IM4f64HDsiuRUh8KWv78Y7Edb6Z
N/Fpfhli5XdY82ZH5ffjHtVmiKoMhC8KpsRKvqFKMWzg6L7ygz64AID/eBcDOFW+NZhPJMC/8eG+
WhDY+9ZrtMHR+5XZ/QKe0qIMmF0eDtjX1xYoB17Ct3TBBmY54RRo7Qoq/JHJs78c/uC08GBqEXq/
AG/UM74Yzl/Aqnxv9n1M9I9rIyOsIeQKEDaPYiRId1nvcd96GjQBwNVHvnWAq/Nb+kdI5abIcgX7
oqWqgn2H123usKsOqCGJDqcrwalFjBULWqH39VJfAQ6raQtkgKWP1YulP49D/M5BkEhHmLqJsE1G
XnoZhcVNvEWzDmmb6/U2GG6vUTcAQgxXZWonrVCF2S3mIghbSCooDTnEFBf81OieWFFunJgpv0YN
arVhNdQX71Yr+QEcWBuTkOArMUdNdN1XrjgALHVGnVp7EORG4AgQr3tGsu794naz9e48nsTmbtvQ
+7TP+aZOGD0GMMOnghkdMSVsJDLpCUcn8Ylc7z2ak3UOauo7whAg9meuLXEh8OopN+l0lNb1c7vd
RmIwwHdUxPWsbk8fXrHoP51QiN97QR3eOnXj+jr54T3gzJ+hcKMo6mn7A2M76lpFOe2b2vGDk6gZ
0FISedsLFm/UTTLds1rZt7xyOC36iU0ljTlSrbR/9qBNQW1slWeE1tQ+/hgPRUFd7O9J4poVd35s
ugqIFaTteDDoq/ZwXh805cpYPupYGYY3crHrD6fTHV5rOic+qQAlwJf7elj4IwASUSpJ/JxzFXm4
TfvEXqYybr9INq+wSk+4PSXbsIVhbjj8/picf+4oo9T3ZyikFKu4aeVePCq4fSGMEFCEAGPDjwLC
DWHVYA09Lp5OjPoN1elrCiI9JCq0EXkRik58ZyKvBZC9i75P2XHbEsXgwXjezcY/L3/qDpOy1tbj
z1687pZmemBMPNhLE+U40OZlYf91M+137yMjtUxAjzHbadSN4VjFTr8Tt5cGFvgx13KU5Jq9Mxk5
ZOdBTTNrRIoSJXGPbAbZMSjBxv2Wew9nNEBXioUctJ5jBS5tu+Q1BC8iYKPm/XAqZF3fChFjVhd8
GYvUPeq4Wizsh7zwZR4UmktlJb93hwlMIDDgYQNaJCcx70aWls9gbVXD5rIhc/8EP3O/rAWGIvHV
8W0kd56Ba3NHoNH8XYFpf2IluBPrQCznEvRuGgLtBtQVFiypkjaNth5HuWn4WaSDx4qlj6idDF7g
pkGuWnXB/pae9DeDAW//QPKW0ue12Tur8YdBuzIrbhqf/09lCzjJ2U/CBG7ciu6UCWY1dnegH+O/
k7tDREcGoLoikDYDqPcrECMHS9KU80aMdMZUhNDtUCcFHghzkH9rudhiKrq6e0svdMn8PuYdLd2H
2kVsW3m1A+WxZ6+J8pRV6gHTkddoGHKTr7007vEVBw4AxoHrCND+3O3aO2Zk8e3cN8u2KdIj382v
zb6ahpy5bBlIRsrpJEwdU//zbF3H9yMAGtYxqDH80PDhyMT7MmFZ2hLTjxEpCrBLofp5oMYxbJ3J
z/+Dq3FAO0d+acz+Vvdwr/QzHEr14P3kwX1AKtb4OciN4aS0vD/w2+P9tnXmhIwKhI2t9sFz2Mh0
RlEL+NRmPUWdpmiRVOyxaEKAYRb9rZ/zDjUxsNPckg6zwznAXOnL33xCrw9NeXEw1pQb/doOG6e1
C3i3y+siUPixQmOCzE+3lOitwCm8qW61IvkTtekXFh1V0BdSU2ccFn2MEJ3jrWDhBS8qZ0xrnaDi
+/ZOaDixL75hPNPE4oE8HGUhwy/4TtMz1XlhjKvyH3vlNILVInF38svfvhpfnR3FjtBHglATPI6C
osEJzJNDI/Xgf6xkzhLbAGZbjpqh9JyZj8sYnQ1dO99pimc52i3VpjQcH0D2wH6urIWrhh6Tma1r
8g4zL7lKGVsW1pn/Qbnr+jOLxV11P3MBao6TrvBYyHZou40u+9vVAlqtLNXJ1q19sM+mySBNbtdP
pLpRKv+yx42UamNWU1D+e6AgbmKZsFWMgiORkKJnPafL7FIZPrP7apJaCuGwf4vqK5/JY5Yw0DCD
ahoguhIpYccVMIB+IYZHrUscF2vMgn3hRAQsXWN4RUvy4cCn3INqu4H/om+p8VZqtSE1/d/o5+Ip
tuAaLXKsjRYkWTRiXhiDpfHO4UQaLcKqTpYcFyzOIPJSKZZamGCMVZ6Np44mYyupUsKP2krST41Y
SRRpCzpfMYE4Q68I1vs1FQ/EDEYtyWx8gca415tpfnnVZCVwqTcAf0mNSl5tsn8ckT3X6/J44bT0
UOcydYsBBRqeoU9At64buGayMnDNamRntu6jS1+4yU6YdFl+t3VAq+lSNWv5127ga1kYlk/fY94/
c+5o9BjFR7tKxpYvXdhIQik+2LtOSf1UvyHR4XyYIcVpEYGvgQ766Cxj+rA1zvcNIn+hnK+Dm+h9
3bxzZJ4nxo2dFWoPHKEgtJG+8Y+5S+dv2vUb8RERJNn5aLoVqQSIfOGT/3xX/wPB5Iwbuq1m2P0R
DHNnE3B929BGDkgTtJ3xirkeZgcIGOCsxiv8iE+699An0Piqm1sOWQlcvagJ8iWjzmGe9oKr6CdH
l+uhQo+g7BNNiSB5U7vW8QvFycGf/gY89nmudOXowMQsaahXxDenWs/KmxOB8tCPzezN1q3MPEwH
3CVKl1gC7L2qZK5sCpfV/padOpl0QPfppzHVMsuzL7pS76GyX2T1vgVnpt/Bu+KKHce8tGeF7/bA
aalqW+GFCJQHWM2e1kw9iKPwIzpXLAVPKML6BA4QmzGqEmsLcgyhO9AOX20YHCjyl9PhfMFpmPnI
+Cjb16W0O7G6Zb7VntBvLxG6dWfGfNO1sayS+1U9NWQUSKvub9BD2IXNYQw8QJDvV24vQEDfonlC
Bwyxaf7vqj/ArbwVD5hmnk1K6bgbeMcbaBEBpmQgAsL5HECqCNjxrHX42XCbfAB3XKCQMcC4XEEV
sHUrCtumSMuvinu1MDn+roD9Cz6SY/eRN83a8ALYFNR2U79Ycupy3kRU4R766pmxXupc1Wq2FFuG
UR6bu7vpvQ7s24JH/VXZ8jvF5SWFOW3831YefJmUvyNAfGaZsWC4/CprbR8QS0gpucUsvqYrzrrd
IY5qJORcx2S0pxTOX7/chjlc+6dr6pbRoqnFXeXZYUjne1/88HiNB1ahGzZyAV8iEXQ8OkquZ9KG
olfqQ1hgrUj5xnegpFnyqBjuJE2KWHgi+qlwIuVj/b3k2svl4tZ+TZklGuDSVu2peEDbMa9SY0ua
4+bcJTJ7UE01MUsnXZ2UxI9h30WELnfbG16I6C6k2riA894ZGQH1K2zXosDqw4mJFBQjajGT7Bot
58uDc6gFpT2iebPd9IBtIxrK869WjW9TNJxs+9BPyD2M0asbT9pZ5ETbBxtWtlXlDVZx8gWPQKI7
2jR/Xfn6nYSCK6W5uNs3TM0c/4XUs7/7NTSVLKUhJgPncaNIdJmsKJNGCDfnyS5ObdAaDPviAl/+
6oaHQf1EA4wRNmqKILYKK+zg5iGNvtU6WlCASe2lnsKtO2XJZiZgwXoJK+SuGD54vHLfEoYEFmCt
MLiUGGjwBZJrgWTNu6Nkc+jVbLrQ0swOdw7MbMHBf1aaitNobh2zngbwATsH8esdlBvtO8CCNWY6
6g4GbCCpSm9yCwDGGMj2FGbgWdrc+FRWlfNoYsqprfe/AobJcErIcY8w/brwqVWrqFGy1gh9OddK
Wu9UufKkYe0I6XPuqd62ir7A1DCzXnw+Tw3XUr5OwYbZ2RTc4BZnZflui3VRE8gEgXwqLUhespdm
XC5VvU+MI+xY4QaFc/5diZOV8GDu7ziXn/+8i8eTe6xSxoiCP3Fvvfm1VWxYjqZARJJN0qI9rxX8
5caXlSVORp9s31DR7RLfX8ESTHjgjOhx1zv44MT8W5vxvEqSf6RJSJLpNBjcCn4Lp86XAWk1/ukG
6R3FaOgQBmysGSZqO79Pv8V1dSoYe1mhmNMMZRRdSZ+tLfmNNLdBeCmOxtso8DzDZHc+X3LUZf7E
Go+LXpXgF1wdE//WGyVFNKCOhDoYFrsv2TUvJSd1OfYZ/J7yOGOjcyjZntuspea4AeRVLMLLOF9j
JIRPOLXrDnQsmebp2nf7cow8D7P10HVm3WZUkq7KRPl+HTUxBL1wdyvbgAnKtErvGSBNg9Kdv9pv
HiHMtnvQanEvmM4SfGuV8awxKLingK66hiWrwlzxSw9khpMdR779GyfqXe2UJmr5GHlE6FzxQrwC
rDVKNv9Dn+lnR/BhyxCjOkUNSnCn4bbvdm+cR0oByv5Kqx8SNoOB0wKIXe1Ff+M9gDFy4G6vpiyE
cKpQGDNoTxQ/33YJ+RPkLVmMqyJYEHp/Yf+PcNsH/fDX+b04tR4sFZul3qGYaCZt7xF8zFLKAnHg
luqnEUfv1tFV5SGsMmhT7zLHSEDyVbDFjqsOtfYbHwk4YOTPXb4w/n73uRnfMRJbDipaihzyRTxI
WXKJ4J/Tc4AYtyhqPa/2946hLqNSzVdwDUkLrBrEadcjyVJ8/k6kImxjStyuH442OZRibenCOQv/
0DvsXboow6LBMA655fXqpNmTengYeTRiCX0PQWy+gXhlyb+nCYPB+hQ9gngwxrQGZyP11HU2cjPh
uhOKf9pR/qn3xA5OitOOn3j0z2G2aPTAQqE3z81+gB8vVGLmt4ZzCLjvsuFqF2hClT98ltn1oKaB
5iHaM67BwSCFQgU3y8ipjQI4uYqypKf912tGF2sdUqbcSh1/O0hL1d58vkgzTYcJ5lskyv+LrF/l
P6bLsktEKhFa+COpLPyboFYpl1n475fNgVlT1aMA7jUBzeewnIbNMl50WoqrbToFZBY2lnHZul70
OcVcU500vwpiCZtHreCPayWLEdOaoPF2trVFCZs4AroI+GDgW1pc1LEr98LauJdWs6hKLtHwSFYY
TQtW783NM8GiJccxOij6sBK8cZ22j4FIz6uSHXyvpTAzWMMxsyzxzch7Df7SjkDSkOYC5QaBjoBX
EQ7M7+YMPLqZLh2nwsJJ8WvtoN/oT3uw343wcAXgtW2JYEW2U3/ZhhLUOExGkwd+9lFtGfD5ySZH
gKgLoKipoqNDeejxt3n3cO1T2vYygIoeI4qnPjdPlmg5r+08ZhY6Lzcj0UDdY0yDDYnRrj67MaWA
5X3RP3J3yNb7rn1eaDhm6lTcVNOfIoKDUI2XDP/NOvPUUc/XXaq9qwTdsZ1ArCduV6C2AdB9lFzW
Epi8MUfUeXBZIJD+U22/Zm8Z5PagwSHkk5Ik+Fxbynn1O5H/DYasVHYyrE7CA9bsyHXvNS3oSHhb
e97Rg5gyLj8xNRHst+zO1Q+/dhcYWsbTy53j1o9guhP4+KdlW4kCwEtJ7HHvYxRf3F+NLuttPp7S
D1QQVJa1JfuSgdjuEgOowXQPgYRgkdVgDbZzaZ7PmCXhIGKFB5DFcou8oriwM8wtTeDOyrBs626K
xZXPYNCAUBmzaz8ELx6vDsGLNSZ6kaiBu24xi06jWYWoehI71sYau6cIc/je7K2wlUHWk82pp8Cg
2xMoZ4O1hGfxVhILRJejQLa7mjz+WvSrEm+oXe43mLz+5NabfKBNz4Pf3IT12qdHMXs09erWNTTC
vRYxOILivJtIikynrjtmG7vGgUEEULAufP1qP3p1CsBOPhPHZ/drA2eF2uR/YuPKKOl+Tuq6YyAa
yLVi3TEAkl1V23EqtMycIh+twRUCOQUB5hQPKsj3EFpPnbY6DQXUEh4dPRxhZGmovZmsZGkw5o3S
hBuBv55rxUiGzs6/r9jTJOMSWDR3dL0vLb1RNPawPEbc8M6a54ggj34Jh1r1CB0naaLWzuK8EX7m
K5fro++P107ZVJr0PR+6y3+bYfQQ7KmVyfjiIvp0XymLQnU5PQEOm9R4v691tZcAdNnCHFTik6+q
ZO3TyLD1HEHf17ooj+UnoL0OTcSqTYAnbCH6P0XKQ1WxrKL04FcqkYTT+w/9HrUQGiU5vAvXPgay
uJaly0nFxPZ4uCDkxsIEIofX+rW+tC/ipZu/q/reqlDSuwa4z61RKzPwW/eKxPbsPnFAfZsze+aq
gyV3BBZc9+p1Dfgf7RJvapQKOLvdcWgNfxa5+v9sHVNtFK2YDn54JK8oI1JFT3wL7vG0Z3v/9O4C
P8Ten9K9TwtTWw69eG0fd/8KGIbvj7+0/Thtd+5ok9jXyqkLNJp6kRcliCWdm/hYiX9x2ZU6JCc8
dJptfjgzJkc0BMxxLPQZeUFPwAC0PZ56eJEZ6uxvkA0B8YbmXj8QJJtynjjyxwWzLf7Yu87Yukyt
r9UpLeG5muaPThK6yBd8DqZWCdcGuviWQ/txqzzh9UBQQ2TsvgJf+kvzAYbnyK0S49an3eEwZl5I
v8h0I6iWAn8tyfp5DUHRiBs/uuWABsIF/MVUgjVJn0aOy38bRszgemwl042e1ZjTMSa9M5eLUAmH
wTHy8ZQFLSS0+F87APzo7hzRkhVHLWLUECsIbA4a+YA4FCV6TGGh9WkaPp5ZFkGtNHQd9gyuBNI/
gAxUSaxJt7/V8vS4iEM3HmlnKKb3t0fO6yySlF80qSL6KWoc9a/tqPUxWgrlsCYi46WZNv+cntLJ
5yf6AzvmsO4cmHmNuAWWBBuXlkH7hmy/MFkOysgDslQnh/NOTCV2NaNl+04YZ5hSyQbXpIuKARlP
ZHfiBcve5tLOxCNW/6VEco7Km5yrK5s1VylretMiDbJ5oX9XlHAPc2TZqNft2SuIKdGqCSrhDsVB
p6FdsezISubxQERYxkBZiQkQ4UxTYVtPlrk8Y3DxpYeVd87sUqfGTI0/ElQ4NUZZwCqTjNeahk7c
acHSIJv32MSvLmonDbsK8Z5RF4nMd2ldPB0KMrnl1RGht8quQsqQ4a+YWhKbW/PkGHwGbiWnbUzW
ExDtumJj28nLPb8etZFtZr+yM8WVizAHqI/jtFofo+N4xIof/0Qy3GUpbLlb7DiEqxvk/bYoFD7D
Ox0wQmLFjd1QjL8vI825uSFK+cWJnJzofk2mbkoUYtzA5wqjqkKQfb3kSNTh8g79CAdDLRmCer7x
TdgcyHRmNnZa7PWGP4Ha3d7jqCSERd0ZbKaqfwIUDgZ9Ia9XguM6YPvqmxdOBrUaoF4Rew55pyKz
tPyDnPPVGdFOvTA9o8jCsquF3aNeKtci0KvRZFs9MHYOadHpLxOcNmCNf8VgemOzlvkfH44ujAak
5xoVzKWd42znhbq78rlmD64nlMzXZPwgUXA0d6HKuZXv83YZhTPjulPTHAytww2Ev2j4UeW5JjMI
9s2AfKwxB+tLZBkSt95gDmy2T0MceF7Lsw1qRorqRNirKOh0TSFs1uwFWJirlb4YFDe6ShvNIsHz
vrsULpwP7wHA5CcuPHrB7JjziAF7l+axSfyC6PMZeLP3uYsLorvw5SQ6g7UbV12+5SdWLTjD0pSa
AwKlKN4OXbBDWu4u+/6TGRoJ9KcYX7Zme3khKS5/wOs6XhISPFE646+Hw9wBfcRIkqcozjMgv2pZ
bKiIfu0HCoEYd8TFLAgEHahnjTJCCTZ7ovzcfjmdUq0OH2Nzr7VDNi1oHoaI6qdJhz8Fftlk/R5Q
KL5oV4XX70hAjZxNHHArbdsXtCLIA3QmirNGM5L6qDggXcUj+ZlpgOpx9DS9wMF7D9zen6k8ysBX
mz5j5YJadYe0UtF35/P6HwYfa1uOfhG28dibauq4eP5LphktdnO/ujcFa1YzgwvuztdfzSm16Kaw
i72fo+a6674HzMI8AZe22MN2EUowZ2XVfPX/aAdoduKWBiLuyPcTlFHV/c9k8CvhCHyMpilXJzTF
sRubghPyC78siymyO7+23xjz8joYRxi5qPdg1R5uQor/dLtvG5RU0+JEjjRzToueZvztYk1DzylF
yvqmpPnvZXp4e/PjzhuBWACw3wosqvlxTrl2Q4IlNcvL4g67rz3CTVyBm9adua4ev9fxJwjXSWTk
uaLM46J/EVI4aa89LbH25l85OYoneJSwXKhMRaHyO5Cjpi9w0Np53OgAT+GiEuhpWI1+0VckcLgG
1Wf04XOtUUAUgmvutydF+dkzz8sF0DqJWyz+iIIAZa0cdyg4itpZQcQvDQiguhY+SHezOpbhy+SY
HTd1C6c5sXOOH121WwgAOlUgN4awN5wEi0zNlDpdoLNg19g5CH41pDf/+uujrai5icz2OICPPZtx
T4qj/btCw5W3Bm/vLNqqg0bI9jvRQ425HrpJPadWKsZ71Ttb4gAuEl/84pTDCRr0ZzTbyPcB7RSL
787/zziTrhec61b2oOyq+PvT+rOEZrXDN1wx4/6fdprWO20w0YRY5lYa9A3CjwCCxjbSKWGMaAHa
RlmwndHx7Lc9n6RPv1T/UJd4JmQNV29z2fma96z7c1KKFZ8gb4ll4u/hF7OLYpwG5E4fAwpg01tc
1fPp3v3J20hK8xzMSsj2vJJsBEcnQeL3ib3jPHLY3JSi/DGm+gpeUoroQfbRP/dsBeoQbQDOo9+B
PjSJ58iaSki0Nz9Fzd9KMfXnPx+ucFtVmAyIz3f+atefVTH7xlfkNj9zWhL66WmyzDtUxvB1wGaD
Dp7eEs5+wyCTtyswgEqlLZWElV0xn8p8W32WX1VPtBNiun84yJn5AXBXThBwepclJj5Vy/pVBb0+
y5HGhTLionRgukCweeq7hsW3NYPH9YQ+xaE4galidd8EtlZQ2078TrHJoYB03Tgp42FMnC11fU5V
xBK0wR9YeIbTRdCSHUuH/WYnj21TgfF56IwUmp40E2pclhCS6iJcWi/UAcpncG+MHGjfKXs0RXV3
FPppbXD0s13k2ApdKxcnP09Mbt0cOQiwlhbyc71RIMPEOqbpeZACGxcaDHB2VNyGnGwPBKu9B8Hr
FLeYHhhHUClF/HiR5DaLiEck89tEivt/uq+qzx714VwUPZZyt2dwxuQ+znytkDDIZLVND8mFcu0v
6XrxA+BgfAkCH+jEwVyd3CYryeZtmV/w3Jc8zDCYKmQ2xgkFYFLJKSw44cW6Zy3rlrA+CGB+yJ9F
PpS2SH9dnuTflZysY94vrXHZ3dQ0oTu4MO6Yq19zMZkSBg3tIdIE0L6kYDC5a5tdILOIa9sEHqm7
L29lST81RGWT+ZORhiUUEPpRq6yd7QX12of+gSJmTxZkpDoYQW3tVgns7k+87iaTjsdL0QXNdiaq
7ejJGR//f/AXKxyLrtzCzvy59W4r+A16WviYZR5OIuLKY4/NyOpxQqhSy1w7QlX1pHdxSCeEybwt
A+t1W+2w7BA7t+5vb1sj1ea2sb1VX0ryXYpNk1sSHGiV8P3Q/8tm3XC5LrnVFzSaptMKn5SirLpY
shF2mTjqzZuSsmuHzafL13EQ1yJNsPw5p4rhAE9uruSK3P5L1DDxMHvO0wjdReWlcK6jwwviSmXJ
4Pjmy3Ei/t/u+F7y+qQ29jwwIF7sk4m7FgC4OaxNb+e+F6GHfKIRRi1y7tHL+9CRSIv3PZPk2IX2
QGNzOjnfBg+jV1fLBuojcJMASAg9GpI9aFTjP01A9cc9/PYnJeryUxawIstEw3Aba47ZlWSIAm1X
ZPQuUVX5cm3eF0e5KdGIrbQeWaGG5ou/fijsSE/mLOnQOj1kLO82ovkx4FX05de0kuyfz+VOoc9r
5jY4KeY0dMHiEq4Uk3cYIRJuXy5Qy5+AVVRgnKy7MBiMrjmwuev9fkHwo38/wgbPGH02Uo6F7AjQ
qodxQDnmRAsV4YU/6zXzVi8vZ7VZ1LOW+p4dweW7w2lvpSFCqXBeNSFH9vCyRd3GZ3KRvB/3fX9h
F9EibpUTUoksUO8RbJhSmeE3SX/NRqBA9oFi/D/lIckmQNcuO9+EpE601uTai4ATihhE9pTn9dHj
73Z0ENOgnUVdIxZHNgR+9OHcpmHQG0l5daSzXdPMBeKBrsHgQ6imdiAJRmNRbv//geaCKqdRtR9N
y9T9fvkoR/2hNIRvUQd/L1vaRCTiRfGyi/eNiTUdw0bH5aszhdXtxNvUnO0mKV8GRtoF7g8cJOGm
4hUlJTJncWtmMkwsd1i9ugpPM3QSzfhKL4nNxv1kZUvKtQsx9KOcsJxRKiyNIDvP974moqwRGLva
UURfAWXYKSGZxnMzAENPLFBoEwAOop+VHgUJkVQinHhQRID511O6L9wOY8gvSqjgd9oabXiQtbau
jq45kRwy2eo3iM3jQSroipYOSwYOOgQCxVlksJCLgE26awlPi3Vjq6vv7T0D8aA8w+T3YKCW0A8A
lDLBh8ynYYSuO8yKho+5DnuuTh+xYGtlS8VYOfY2w0UOHT0s4qUhOBVeRCgLeh3hggctkxEtpcxS
d+YAgLawTcAEuHOf9IwVzW4DGoxS7+k3urLOFMoJT5nUSNCWBZtnar4vQNOPQA8pAZjXqBOprdZU
+x1Tu8nXv0uoSosXGtkCgZQfRy9xrRR8k3BeaCYV+CcvoxbymlZYLSDJRpGdZV1d8HOqMyrM1DpY
JaK8wCVUCgugUhSPSTG1kS3U3rT1CzNwyQz0V++JP50ewdYda2ZqVjdf1yI5MR+CCeXilz4Z9rKB
06YciI3/4AjQSrTIJr6JngHmn6rLWidA2aPnRChZpzBNF4G1upH4piQ8THUHwBUsPog/0E4XB8QP
xEtvqVXLUEYFcX6a5Nr9MNhq9gx3fSAbjjRpPXFq1a9wxznQ4SP6WQv6ZAqWgxpo+gHMxSfD/dKE
iHYEHuTVdngg9zUNVPX6O0WYTcr6lcgJFbjApQDKpO+4S8RUsZSQUV4QHSuCEZ5tjQzPTarCWFG+
g01PYHiUPjdxpUXuubHmLLvXRWkwTVEmHi1oXuZqoOSn3ud+h2yR8cgHS3rqhkNkWdwdTynTbstt
GbrRb/df5TX1or02UViQ2B2SPt42ykRebRCw5iBiSoeGQnobSPpn9w+xbEP/O775p2qG0+WDbR4l
NEGFp/DkMwURCAfp1O7i8ls/OY+WJ+Fx91vW4pY2QQzp8KGz5D63KMea4/x7vIs8ZQKu3pSzuOMp
WP567rZeVboSoB4OVjnhfz7GhY1C2frAm5eyf4Wv/JiFxpWnQQ8vCWLZRrQr6UIUUTpGtHlKqqs3
HJWWQ5B60adm8zGFaV67lnq19l/9eP7q1liJEOx5HHggt8RWoxlaKI7PCpVpPjpOaKCchTdI1F1K
XVJNbHBnqQoSQ7pXfGV420lGJf5LvuQ56gJo0pB+yVpn72spz4sQhA68eyc8MHSnBG7uupE6Gr+0
g31z+tUhK56RRuVsa9h5vxLbSmdCHoZsq3nQTxno7stERuh4ObbqRzSlXINVzV0TRq0H2OvwICqJ
xYAw73W/jnRbfE2FWLRfXPlVlcmPgzr7nNGOFsiXZG3qt8raoltmxzCd+SkKb8tngtB4vJvb1feY
aGaljmWkJssrvexpNQqvXRh3wtcIBZGjfljsnycr6ZypydwSyDVQeivxRVbAIwKkphW/ZrpXd+hl
+9NAACZ/Wn1Snlp8gQW5HQPTLThUdyfjxnKGwuxEGVjhyuPZrRGe9C2xeHVwynDd5AKuxA6wXRlJ
H+PD8ZSH5NIb5iJvnuPwWmTlU83nTPvJnUbZGHsIDjyIo0swMAuw67E7/oOOiBSV291ZjItiTC+7
kDxO9I/zvcIartlv5ucQQPemw3DjCmLq0hH2X5fj9ej/xN92VEaQSJjQNHeAelK+s7/KtB+HReL8
S2oBhGpDeqficSXBwBuoQ4SNgUrqwskjc/rIgfFYwloL0kxWN9WhrtKePZDE8iHPwiOig807iU4R
bcMrpWJ2qtvaDsBzqjnpo6G3/whior/5E8fgguHtrBP40FOpHe6cN78eDEd+EceGWudMPp9NlKrV
eFYXbdglMOcg0S/qCOiyMGDhhFIr6R/WT6w1VpENGpBqvLRsr98/X5L18W6K0XOjNkY1r7cUXaZC
f1A7Hvwaka0y5xMrWCDKM7ctsMIU7Kx5/MhcanWpVFWlHo5HTV/Yg70UvnygcPN9zKu8arWjx96e
ZAqZXscXvCyDQtshNV5L61hsxjCQ7dQGi7jFl2F/yJ8vZt/KzJYAlil5EoLtFnac3OOiwFdKklvk
TFbdNOBRaKP9vQNDQdNAGzN71FmEipPVAwlbw0UnBnjWPRIzd4K/OJffW8VbYFkAu/gtb9p8LXSF
Kd8DS9El2yKEScTUjL5BIO5hVGnSVnCGDLTBhOgq03DatVOgJHZ7+ZfPwLeADnLeaP5LY1qEYmrD
gt1VMPfsRMUpTTVAvdnDgwk9F4t9+51j5CuHpMPWCcoYjGtJPVGt+0WKNsWjKTY10NUaDufcSsIa
lITHwvf6jGPlqHZFozsQB5B9SIGES+RUKkkQuTS8laliAlWB7ilPfXtnuMupij7BrbExhsU6Hnge
kILWa30fDLOG7BVOptQAbf5msudJBoIATWzTW0969HOrr+NAmDSAsuGwOJ//zC4efj64IR15CDdZ
qkqeiFkhoS2oqPP3F/JLKGjfkhfcBAyXJCBYY+uD/IP4TMdSFbJu9ruvh/5OfZnnAMODzZDoTTGO
0ezyQOxij2tMx+ICw6J5VEhHE+Em7hP663T38MVzFjUxInYfkEqbDvfusuvMOvKDuKTYLVhJezQF
fAXeMB74zwlvgwiQiTppV/9p2DmWsVhUTqHEjZyXM++uXn8Gxh+wMmSyFKZZMkgXSprIj4zbdAOj
lBndjB9uWzvEKkqHzjWzvlYwPbqtA1Bd09VJpzuQXLNBuLdot341ektJ0QprXZDsbWMykq6FrkzN
MtSoj+7DlKiTC95RVPBGj4vXIcsj60qtxQPc+p/ivu0t81KSVZKZDV70TEJPeOdMhGY1X/ZbZXKq
0m3WnjpkW1ByHdG/Xr3lGgvaUx2F2o1vr3h43EqDUNbkGWfiXmpyS1mt/BG0nS3NUW0oEXN5isTi
ZKwki6JlR4kuSC7eAiZDl9zLJ68yEgolgTI9633DdVSQhRfIOuyClfjFkfiHOP9uSRy4MaIvbu5r
TJO9UPi0t5JEG+nHizGCJKUt34rqviD9JHb6XhafItqfOkRVqKvldEVisz4nAsvyAVNplKdQyAtl
p+A1TMWKK5yzh8UohfQaRBwyuckk9Y63qaXzpiWIcHwPtlW6+voGotqsqOQPQzwjAgtVkZwhkVlq
dWHJCEHpSIPIPS5EdKSKosAgbF+bTMZ9rtfKKplMXfcHEpwfqC8opei4PwEqQ6nNRDI1TSD7cj6M
Tv6X5qnrFNKBEjlFFYG/MzBr/bxKFDi2jWxjW9OPNGXTgQ6JeW8vtEi/rJ0UfifOxJ1DXfuW0/w5
iRYSFzP0gek3Iyh8U3d2FUh4JwIrhI/2PsuB2WUI29QPdszHiVOeJEA95q5o/5Ui2qZjt8QS+dum
xHAU4t76cFdHEY985GxuaVt3zXOUHv80JhJ/NB8I2v8XDsDaNXN+fJVyCfDJS3lUlZV6q5Wckqpa
PEgnaDLwsiJUNhpnejNW7zIOwf3WKv2F8yDE4Df2r0FLvKcTndKNIEuaFgEUoNRaCasYCqvCTGhe
/uqPKFP7C//NvtIJ4ZUUyAuxeXh1ZnP2QtvLbRjsepHCCCXTuDHt7fURYNlCAxVKMC7WnKtqAldC
BtQqhLZmfkcdxmNZzE5vFwo2ZvvKgl0ufoIaIF1fVRFtGsisnWWCKm/f4AduV+x/xeFY31m7GkzU
zfymJ2hfBW3SVgZBpnJznaTGgQ8p6QsXs6dU3c2c+e7vtvDuXB/jTjHaR1MIRDgRC7Gu2YXsDZG5
ww6MQM7nxHVyKz+i3euVhx8J4MsZUy6fyMWrfOSoNyU/F5UGcxcCzvn/accxeQENGgqcd0c7Z28L
/lO34CoY1dnXU0jGriAJY87roEF0vSoyphiv863qj8t4cv0YsHcITRU/VcGHpEJiKk5gfPMYHHqH
LMvCCQCjhnnIe3WY00anrJd+Bue1CMpnPu2dRotyfyhzucJ8C+sGXc9BkYlCIKFC+OcmcmCulGRC
A5Cy+qpSZebd6jRnv5IJjlhpTFpgPbX9LIOZm9HWtYbbv9nTuwvlJCjEOvtE0Peau8RuAW3wBo82
nsPpHBJr8U9sK4hfEtQJrqYbLieQ4zCgASQblt+P40tdqadXeRqc1Oe3nBZpDvDYQ7AqMQBg/PRl
qyQLrSlrHNbHGD4MfalG7Dy7YSTDcpm5zvXYg6gDHnsZDMC3UhSJ/9NNmZ/agFWdu/kw4wVMWqEA
URLkDKZuyS/nLkDKw6IyVSy8CG7SrtolojYjWubzWSur4z8Yk4mTjumEPKuK/oUZyEwr5GtVB62t
4V1OcmQpGajG27EkHIEOqq0t3ViUBqSoAGREfJE/zxRr/O8xTwS65keJojI63ZKU95laDVtCuAUZ
hSyfkOPOhocezCHxuSm3OqfGODHJQr8IDek/ZtDyD8YNdGJ5a4FE22+F2IYQOZCrDUHqZo8AVh9w
KNzMonxC/oJ/smmBvjBwLjHe55WEUMiyBi+7+VBpS013Arq7M/BsZ+fVteYcA6EBSyGlSxfv2cSE
vbVAFqVgUh2G0y3LOzWPo+1MQKQQq1YZhimPEeYxT6ndeB77T/RWgud3Ty3ekMDlg5ksbAYar66h
QPyvyDWcLL1XQ/7Feyz/ehhymcPsBPES32f+hvrk4d1E6Q88o92Nlw7pfc7+BMzKwE/KUXGLRb1d
0j7ohM5mX7hRirODRQZEwJupWqBZJsHL0OCcx4XGEsGJq4OHLF4PVfV2LDvG0GepPWF3WRbVT2fR
xtaKClB37D6YcewCgqcAOy8Uw0JW2LmWc9frLU5ZH+Lja/vU49f4yv9mVZN6QzsXITdC817mfati
pkQRHefOwCHJFOPfHVZScfH/2jyAv50q60kgYu41i9Ie8eXWuoj3jb7+UaKYWJJp9O4uew+Jui/M
4Hn5kUIc5WGTAjhb5VILgw6ngNzt9cNGdSx07iENFsZZIv7YCfg+YxTCvWBDIduQu0IiCOQDn5Sz
QFCVCUCTHLz5lJUpb22zQTSiTnZS7jSJ0lM7fwjVR8KFrxf60gtQN9iy89zqaoWengHy2gVmsbO6
NIWNbr+eTNyUzO7IMPb7B3vdrAtIXfsJgvGO3+aRCSNlYAk12iRzoR85sJ2cQ8BaBkckQToxzasQ
gqb10A8oJwAbJUb9JsbTFfKNyuWbBs2B8iO7ByeH1q1M3D6YrShECU7aDlUMovwURpenUItKmu19
xP5x9UFUz+9ppyy443tubLu6ioOA90Q7ZQxZImpRQQiXlwofdD87tUueYKMqQ7Js7FfvFAGzK1zV
J6PnZSD38wRyMcUs47ho1DhN2EvAOJqc8vmzd8+lDiPuTJjDNNJaY5XNcQiiMWnXcY1ggef8Pdbt
kwyLkeU7jomc6R2opAWBYPvMyr67HrGl/OLbaX1q7ODhiD5YGQXwau66EKAnU1VZXGbjVPuYo/Y7
DVkOpfda9qoWLl/6zdaCtTqBH2edCZr1lPMUZNZK6b9RW+FFmZDpJ5JRkO/O4ZZ30iWXofEXZB9F
DY5gsDLxzWyIKnPKZukIoO2t1pWpfVf6hFMdPRrA/1hQK22EDs3AYJwlfBsO4WED8LGdC7lF/751
W9GVrSDG7m8UetxjqKFzqFq0+K9VN08WKBDJTvxSdlT3Yw83/Xp2oiygBnaHkGZqsgJv7V5Pzbyh
W13NIQUcgJuWOs1LcVh4qc7ElvnaRqsL5kvTRnbv9yn/G2+wjJwNfxZo/nirTUJ2z8srRNiQRfUI
b84tifb79cKym++iY686/YhNie+rAeA6GDQgDTmlFSgsw/syT6zX82zryf3pBhQ6GpMtpTRdXJn2
5/WqS6k5R2skl3TFYfyDSgSbE2z7KSNPY0s9NCT5lyOvx8yGsJOhIxVYJsFrbb8fstNeamw/y4a0
Ww1CbhGp71hNloxbX43afp9SqwigMihycXJNAopI1awc1bQxq5IbLdEQq81A07nCkx0StTt0X3q/
LOZTecsstWaeE8KMO2HHrQDaLQolOBbEenWCH2mJjTvfHBn0mWvXHTRwL7y2hSGb0ykHreNFRyBr
E8Y0ZmAYnvwiocASOCXF/qoAeLs//1D8m/PK70izYtxg+qhRq5VJrl2IIPq6olbSJA0L6fzQfKp1
F+1V/9p3t1+nSSBM4u1VbV/qsQgkLV4hh3x98Egq4wBAxD0naVKEQYjmUfRR2HymcZIPOURCS1Hp
zBZeJMc3Iv53cXKMelMM5IC0cBz3Z6vcUTTpRozyAEKoSyjn3m6Be86kobCWyJ7Hn41iFeSMy+HM
c0Shsje/e3ia6Qu8IX/oGxbeXR5CWoI/4i8UsGgxZPQWFLCT4tqIDfTu6NVMSPkVOb5q7hm6ZnpN
RsJb6rSGM625smSTAjuelaEJfXu/+0OZkhfQdZYlIU3vqH5fRP558q0jXTG1KwNoa7w6YpNnmxjU
UCl6VFZke5y0z8gvOw857GXqhJbPG+jSrFKA240yQPa86xjGaFNGl8aYDI3zbVd/ubiivsr5TMeB
d1rKWyJwIAh5qL8+UGgTOdwFVETOAl/Y9wPh7pdsq3KYznTI3iPxHQb8aO+CkMNWQsHSc5pw732K
ENGLkJGzGER/IbSEph20y6JA99H1DcXF6Km11nXlDN7hs6UnCiNUHLlaUCrNI7BbjP/qBnG0thhC
FAz1H6eBgp/M3p8cgNtuSgdJxYBq5hk67HF0XLoTWOA1g0Iig7qHkBO5R3RzzEfUv3B81eV9+WnB
yoJMtqdYT7XrW5MZ51xAmZVSqUgKh+YViTP0SwSYzkSgr+fkEzXBOzhBloQXGRf/D5aWJ5Yi5r5z
h+Zf1SbnUD1gMx6NorqOg63KziPPU8X7qwHQCH7u9Cr4lsrwZAlpVAd1Y7wT6KVOynnwisun2j8y
9fn2KqJqMdxPun+e8FX7S/Acr9cvsgHQPznBqQVj0vYb5ILTp1SEWNHXZVCjgFagh8VqDAIvtngw
34Ihyualz5izwFDKGKJAwBJVswB87DgM7q9YFkA5k/iUImPKp0FCyY8oP7pG83BSwhr/j//X3I/C
RI4zQ2ylOX5sleYISoA/CfSNwrKyfcVBwDnZXD0Hoce5EBr9ZSURZsrro9VIvkJaNFaMzGXtcB9X
WRbQir7ZtdwiuONaJ6L0bVN4DgKv6cu63Yji/ZtOqyw0Tkrkg68pnjsBUuaZF6qZTT1rshMdXwUw
gZi+ApSuAEUYuoEsmdfnKDvCHryahfPdJxhJbuLXupVqRD2eQrfrQ3xYnap83f5CcSx2T8X2+ZxK
fBMQKcxZ6I7/bjoZ7V73uEUZrJ3thg5B913FnRRfEj1yWuSXu1I5UjtcqZs6fmSS6upleMvc6bsz
pJbdwS44teq8ne3TAxSFly97Boxi1yLoXJD/uhGJlTPNh2NsIGq/TunIW7hugn8cLURWdwF5Ktre
lA3d8Ck+x4ELoajmVUQFHP0XaAcCsKB6ejfXhlhRrBxnVUFBOkX3kROZh3if5sneppH+poJakY0l
nKJRihj064OUd4YRBtp2XIVt0h163P9L3+goJKBXVW5jPMKeeeQonfyuX0jUcSTXQONghl0yK7P0
MDkyVojmPtOK8K4fpO9uS2Y6shIoE+ixONz4jebjHMDTKOVjNBFc8/wJI1WVB7njrcyUQsKtL5RS
OQ9Djt227mJ2Ybwd2Vr4qO95qZNEGiRJufeJ+HeuiWFHiQfVoFKO19K98HhJ3mPwolKTRWckJvjT
MwZYAfoNHaFMV/FJkcki8MWXboTgF9TN72l8aDulua0TkKncWYxk07k6txQ1Rgl96lm8lBZTbX+D
47AbMiMPiE5yG1x54UW4kNrVLJ8m+B+4D+6H1+GJjknjzWxVhVuXNhQkb9Ta7za8AuGHvVZ5T74y
CyCL6Srud+64WUkhTUikXFQIaTKMy5YjFkKkCo3PH9spLMTu9Q/IH7hgEASoLtIsBxOPGFfvmLiJ
Y+DzCH1U1BtgV5Hnh6OUxz/K5LUsAPCNNOoSoQbo2r6F+jpx0LG9SrEZByvd4eEQZUnpCBK/GHxm
XRNtUoz8gyQ+zs74aQeWSKhx2Ix9sBmp0zJesESZiIzH1fbLqgANM4C7v8GOnee6ob0DZs3plNDM
TO+fW0B55OFjrTKP6exQ4FPhI3YPIu0NMEedzbstT/A8u2ykSl12kvII79P23Vnp6+lgp6xnAx0S
y9YcbVq4eUca+bGE66yA4r2pXU4Vx4X0T4pUWZuhQT17Eg5axHXt+burpTtBF9QSkGMqsfqxaRv7
K5Gy5dYkQ/bEuhqvp/tCR8rQ2FaAzaYnfGK+TE5pNKZOPQThKIUOjssvfpL4gSquYiGVNCcdVXGq
Ia67DZRrZj+hshHxtrgzwKk6tUSRGp3wpjuTPyVMJJFQ02hlYrLlvOyJd2FeNs5SEA3JyiGuyBPp
Rlb/xp4L5JNyHwdGg2LJAEmo0QXN/fInTtahmS36tfeUDV8h4Sms2gsx/tHogpu3L4Nu1YqRJuUO
PcQtyS8ieQ+b0lgfJrLCykfnRRy0qrH12bbrC6kCG+NMmddwC8QDReJ0cRbSYrzKDFQEP0QnXKWN
61HZshd+2QEv/vCVnGSJRKmNhCZriKrJiY1Xyj0+uJe2dwMMGBkpIBugBSY1S/nxIkNPJua0GCEQ
SMTRmhPKJw/yKITTUzfeHRVntAsWkiJmRJ2uBhrssdNcLSZ+ZL21X9AO7KE3wTLO/oAWol3zQ3Sp
JIs5EseDbudqyd97NGX9DEHVSG1VZCyqHRfPBaI3rFLlNdN8qLrvYMHf9dbNKV/YkLUTIQWyn1IG
LCpFTyEIEbOOjG3fyZ4mxv8FmQJzpq3YeX/lfkqIh8OGvulpvYNHnlyj0b5YXwPTBszKIz3TVjr9
gfYDJyafaZvI9ykKB6POD+Xt9uMoukHg/AArfUwRatIavoorCNNtwBRR7DDhMTHuVnKumS/qRkRz
JI3nEfyFuqIell5YmeaGgVbwCqkzKg8XB8FVgERYbAt0YLbx9XxP3qBTPCueiU7/msTd779NpDWX
PigKCr65aY1oM5Qll/mvFCGS/9aGZogop6hqM+zHpm7tEagHyNHtWoEdw7seIQB1R8DomYh+Nemr
zT2JHJSplMfUtx29ZxxXCI5IXmzHVo9YKDEoPLvTGQdnQW3hk9T0djUdSN94GXhjH7AQMe5vnKun
HWCNVUreX0/hubSuBgjRnE4i2Yky8LVtqrAsdR9bli3FeqUl3i1SJ8wj0bx41XERWnNcxdoYIbym
xW4IfI91Ow1LPyjQnM56pbDem6JE4dCXUpf5wAqQa+oWnZzNDXhk+YK42CstemSFdlo67TyZx8tO
PG2xKcW3Kw9QOT/lD68mUKY0gPlQkbJi0OpKm8mEKfDLgBxDA7P5LuvHcURLtJbCqtjGPQO8+6wk
bqQKoGImUc6zz7w929Y6vP7QgLEP3sgSh+K9JnaThRU4c1pAg3F6jPMZG+dk4upVtJgmdwvHeuYL
sxA1wpZ+eT3fFwIZG93LwZNw1+j0Qc0YGgYlqBWGYJYjHgJrMI2HosCBcfrCqsyOATs4BEBEOqJI
0tLNzGWz3RjPlIWh6ts9Pnl3Su42mC/AIbjT0lnXDjLzVK/feXlpTcyY/g30929YT8JrIOFwfXJ9
JX7qdDNUjQuzxM8oOKs1uwuC+8iY86H0NDGTmXVXExakxSeoyite3qRnGPfjP/8QWUCbi6VVOKEO
e9f/ayxm32/y3kSQV2o4jbczQ2AqQPvJidX41K+EuN0urXbuFGbGR5+MO9FvLZrw3xMOryTCOhto
xZT+ujjC5rS0jmx5riTq6A851m0alWJ4lsJvTjYLoFmmFkKGc/s5vupCn5Nhepsa3L9uzzexxf7e
G2jtxU/MuTQJiG1/GJW7RvWeOEahWuohHKqYl+EzTVadsLZQXhr35q/ZiBqyS/S1eQpROpllgJxB
FdKq4MIn9WgmGl3awhI5IHC/ya3+lU5yyT2ayAoLK6vz2b+W2sp8xaiJcfCKnjTx6hnmCCRywUM6
jbTZIQq8WeD5I7VFP583XnKT3Ob871fTn1LqmpEvLMGvExtD1zxtwWgYpbl/ynvZRxGUiE5UNuhd
mBtwSLX7eMI45wS1cyUoGrd4zCCPNIx1EUL5oTOK62ln9cFld3fImzGYIucZ/gD+F71U0q85/nJP
EgJSREAgC/CZncbd2AzubAiHcFnT6vcdH2OtBl/FJgIBXonBS9SbUuAGOgvwPzeUsBVKSd8P5vHN
atOyvL7MUVudP+QQdXE7EpTPGdYqEBhlBp0GshkY2l48XBlj9oYY1WOLUFw+0FyWWA1w1sQASqpv
abQStUE432gS5uDB/oZq3OJgHEWZWleUqAApbJ9b2TmSy/5quzpLsJ381oIwdYrU5T3rc6KYyUx1
hk1ZxBFt5tYrcCuF7VjGoCvAoy47jtu08l5Im9/rXafhx90Jn9NfcvMohvaGju91sxWN+CmMvuCx
ck8dujIGjRu3DwoL9O3jL4CF/oReyOsFAWAVVv2QKZcDIscrengvcRjwnjmKtQc/x5nnO3eCG/ob
IQOxit4T6DFWfzVtpteUtHtJ4KODmsrMNf5yeGrS1qQiZCwst06l42Tqis8WHWEk/8FLW37lubTf
k12CQaDr0Zc4l71IxMBh7BGAC1eZqHtMK62JfqoFniRks8404xZOyoxO+anlOQFPE44NvA8ASDRp
3occIXJvAbHauxEhQfnSmTL1qDArCmyVMgHLTfYNlm9XKvcNg7JX53eLuuQ2067fvEmUyUtnWaz9
IKnCil5ZXrli6MtnvEHdjD6FVm+dAxfUbT6ExjA6vGmdpaC85MUn450494q7hfOXDJ16FfOafDS5
mXBr+gNtNPXEfpo434VuIMQh5zIDwFmXA/TOrpf8BeE3zdwaBlFDDchOLTuwHCaiA7vFihWKqDQD
ONM5FckLg+abFWRS9PsRq7RUiTvzKos5J75QH7c8XhrQuiK9Ai6wc38JFC2s4gPDYPDBs5JtmaIl
IH38V/YJrTc1VULpn1caBt7agMKQFectEbARML+Tej56I9ewLwkzevrI7ZbHmjxyD09HwLfPbPEM
TN3MBFrya7oKl5byRvcPKzONiw7B7WbO7h+myiA9thQEoKLga4kxc1UaKV1dMTGKeM4hY8EQ0jQb
T6j49BGueVq+NgM5pcsauGSqPdk74q2GOD1c+2cFr3zefxzgRrsGpJS1BmPFHB5F8RjTnl9aDRsQ
uY+EQ7MUzAW3Udl/YEyIkiORs0XPVuIjk6hWdyK66cRls11dDLQeSQqptoCQ0qqxNnV+Y1PunZOi
g1gPIJ/1zsfLSf9FFxQ4lVs4g8Oe8IsPUk9syDn6ALB3TKgMcNRXCai0P5MdLtv/wcspPJ0YxG9l
7AVIvH298srEyAWzC1hrdpTQwgqpiVKhwa4N1tAuagKMwXG6Py18jOMFny8RHJR68KT5rVf+rbrW
XPxfo0vxUKI8B5iGs57UhtOsUM77nC0Xj0MAhLkMDrd5JNdqmr2OtFu/ggs0nBnptSNSZI1gkQ7K
NcFOdZOwdMGdfL9FsFhWseKKLj4+JPVRIKMXhV18C5G8IBz820zIrSGBjwuLYHpm+oPc+y2zGDnF
Rmb/p+Sw5P7nf8OEMULDKJOvv09rWtMh103K2qXCjgeU6Vi/NxQ4oQ6s5/NteTDPp/7BpttGzwmj
bqq/nPa1KACXNdjP45ilVOaB4DDkANHksOAumNBFcDoYi4gRjUiHf0Dv8wVVo0Vp0cgamE+TW6V8
A11IQmyFmz+PhNw0RNRbK8auZPOswELAA10YvwETxYk1Bn2sssaHFaLcMhtlOaWEpOQBgX60cBVL
CnFva6VM7vo03IlWqMf01cTs8ZyrZiXCFNVTx7UhzAbVQPbIgklY/NOMUBDxMcWEU3CVNNnm6SPd
1VIhZ/platrBDGAscEZcb67SComLoYkWlKQ72IXeQ9Jwb67/KLajBiJEGdklFjOOuPm95Gx3Q6iL
6rLqgaVaMpWD6SoqHnnuueLMjt3vF6Ruh5PYCFDwpIRt4nztq/DrtiEpZLHaQPtCG2+x8/oUWBfQ
a9e3d7xNHYgF9/8rPgQ61ZY9RShXWrvzY4oFIEtqY15cqMzrWo+q1UjulmhfkXf3Qa4MfMPWgXLB
V8bfl3DDNXs+IBGOwe7jT2+zUaj5UNjvC1SMBR+1sAktRtPOP8v+34k74B8xKi8ks5HRVNL9Xh0W
/4IBq6ubWnFYjcwWulc5PljXJbSiXCkhd9XL7PBTpfd5b4nsAIq7lJid+Zt3kIanH+HYOlB9677p
s0vYfU/wHa4meh5KSBMYckN1mSeLJBxHPQ4p4E4LLM44g81cYapb+zCnTr1AMkpQJZJTwi+q8aeT
J8nnbgpujNkuZrT3f2iX6ukRDiA/qxpGN81t38z1+zElCG9H8ICFocE/U61Wbbevec+TLpdV6daa
1YQf3yEOmsFkLWXQyNKQhm+xmn1PrpyvDDRXvzxezz8F1pdzEUv6dT/deBN92qz/tNq3RMQa68i1
NLurN6wGGidND9mOQJDLKXjHLlPuU8Wtredeee88eDbrVKWeTdRjgcEGJwY22F0Fr0wrY81oIxx9
kF7KrKjHPz3wTlGDpHydjm+A5DtjbaU9V6a1GmT6gmZ2AE55ROOvjmC6DUsUw3cGjAdd4YVi6MC+
fxzBieajW5IRCAXFhYIKTFMmQ35EaUAak4yN1PBVboeCcq87F1OxBcu1LYsQDmKO3CczwnSv1a4F
Hthj6XOaUWZbJZ5bHa1+9302CPnoCxR/8cUWgNDiZTR1edT5VDbisq9fDiYnR5b1N6di9JX5idZz
XwL8YHK1GyTpz84pYyUZBf/9j1hn0P/YEaCjHiUDYR0F4Mg6NtZe04LgMfsobmsDUt/i+JjwPgHx
KqbLEITQ+9Yq2HuxuUhKOV/9Ovwb28SrJLOsWR4LUPWmjyPjYsB0UJhmWaz/DVMv8++fQOg56JCR
TtJW4h7hV7OdneTKWVKu42JsZWqZEqO0yRsWJE7vjidrerG45s99+Wvx6bFmkChV/apgbo+dwLa+
tXUQ8A/OGC6oM5j7RW3cGFe9pGCDskmhQzXIurmpNvmbM7djMgwatXBiyOptj6OIkKcoq3eI5fgO
gXZXpM/+yxud8u2YPxvOvYdlktOqJi217+ozpDSxSC622UjP3xs5r2A/z4l0akffo1JRwuAsr8wY
eN7nlHjcXXxI2C3rWwK0AMdTgww3vWD00QSYjvv8H+Ar7Qe1CbqZXhyA4OcQ2WXWJ9gUyBTaGywC
g58C5cjGDv2eemsJQurUUTMslPuHtMU7imS6CAPH9sokVbV0cLnPJtBlMSEFjdQ7wwWZnvsk8QUq
uuaGW2GyGD0gIr5EyJ7RA9egZJDulXX+wtGyh2A44/8y8Pm2xh2pKU9lFeJMEzh67kVtlpGyA37Q
14drAyyR+rTrLgpAUz4z3+WtN0h3P4ckUX1Usx6pFvD8aWoAnuOZsgDwm+kAYDG0Yeb+dQRl06Eu
IPLLOfig0LeUgP7vWoM3Kyqde6ObBA3KVxu09/0Ki/tL8OfCo08BHQOI0FoCrQODzZufzQe5htSP
2zStKBVOejMjJfyu/uQsu2HRKoQ1ImiC3G2OaieVqNF3O81Zvkme03huYOUtbKFAC0sLRXIgkDPa
R7GWpy6qa+h2PsODWExicLmzQb7Zp7feJYMucEWH/dRyLKxP+y3td1VhdF6hEAmAKbxBkjk4Wpnz
C3hG79SDLfvTI3E8+tXu/qsWd0J7T8FqnRitPBpGJEuiDErwQhkb+Cd3dYdbWUDs3IJn7pltnI0k
hriLHSkT3jo1U0Eu08MMBH97PXJ9t4s0ztHjQ5PrNQ+4nfofBfqfeLjK9UVCo+8LgMneuqtftmft
keWzlQ7W/bu122TNQFGAhAvi2x7ZPx+36/nbczNRMVYvDf9bjvH1vqXVKUEUFFeCfujdIXAGT5tv
hVF0gLpKZQmwfw3eTiT6V2p6HqLgExC1gQdoX3Bi7AvKKJFmiW00PpQa1PmfHkSgey9Kv0fq9NbA
juWUVQNd7zRcyt6r0SfEfFVXYentUZEdkGzkB/doP6pJ5hkiswS7DXESDOe9lObjJ6CMixKp3/nQ
AUV7GGemeW4GkmHQvP425lQYdrfnc/e6f4UsnL2UhhzAxqJJFdg4RkmNhv008UW61+eCsPHAuFaI
u3NdUTWYaa3T3VDLNcAiFtuge6+eVP60LrNMykXqFRVSceV7RRCAxdVmnRyLxheQu+EkLVbA2YcT
JTc1O8bcVU8f5JtRRsTHYY+uVnBkksLr+xWhP0R2n1MPl04Vm2QntTtjeZAEGCqIq0qM1RYKwVEh
p4icXRI/mcAZC75Y1ls069p7TiNrod0R6xE7mkGqIQ5U3lkS5hXkmcDh0hQvJvCdKmc38tDvyBWp
3Nrn//+5hetEyl+CTMsvvAWzYuir9lh58PKrs0yY0Uof/W4xhuaLub1LrpUFtu1BGV29sIkQQOob
U6TcYxBXD5qC1aZQuA8L8KJukvLmWdZs475WvSbqlqQEsIV6V11rumkazUXTWqHafVLLt3sqZhMT
JYydNZ+6cLC16u5wS/IbXBDu3e6T6WqFH+ZvMhbr7emz+NhhvMBLh72Zh3NtyzHjEqZRfkNcMszX
gxUoHg0VyRFfCdPshGPnY7RTbZphdWnivZUJy/b4Zte7d1K+IaGRl8I9Il/UB9Ao8vGfoLdN7lU+
2YKKa3CcHR1DlAAQkHjQzHCV/wo7z97YAUg+MYXoh2ICDsSzjCjBq30yki6QgqQ6x4N1fTYVEkcY
TjE94HD8Hm5tP/ZeJ62Bn3w+FFKuBwZ0qhEMuLWFucF5Nyt/qes4zumwcGSmNNnCuVKxYI15cijK
6tGsRgR+BWPBqZM13FnR2MhU/nHAQ7FNoD9nwMK/fmIx1vlzK99cdUXNp0RVAqgLAWE7A6hwIQXG
jL0anbojy+gZMCf1xCC+47TESJmacwrqxQw7UVq8xVDWJe0Tq9MeQArC72/Up5JHjF1sawnNyW40
BgK5xMZ/6SgC7L6wAwubxRLkYqibZ/UpKpCT36dqIDxIa9/d3ii3T9HgJGReR+NgDDgFktiOLPpo
JoG7sPnrOf7lCOWpZtNhoW2irxYlKDrc0cfKqZNKjzGpbLTjsi5eDSAWlt/B9uGcXaNtJJMMJMJj
0jD/yoOVlQayC1maSQO2vMk7OZlHc2fW0QfBszVjvVgqu1qylm6VGJ2Sc9yftC1P/GiNGWg+oj4M
DZFl7oBe+ckZETW8QdciSQafHb0MGV8Zw344OJcg0bperYrRLm1IgUhNYDV0KDF/Kk0+vTNcIHfb
tZsbL+wz1iANxMMfM3AM38hSIpiRRKTQu5Sx/FpV4UhdokeJQuMqcL7SOA5buKyavSF7XFnbsd7V
UVTERA61wXs8uCqicV5F2rXZ6oH+EDafI+VBdS5Su87bi5e2ZkyukSfpX/UrrHaJBgkJI2t1KByz
yNtmk4kSCuJ3uOhc5p0Q61bRQZoSf90vRLLAIopgW8jKMxpRbzqv2Oy7VdoRvqBBYwxstCZIe9RO
TXfuZjX1+y1oKoKr+nljaCjmCFIjwM6Ya+KOc1DhW5ikr1s63Zpp3XBl4Fi6TTUZThUTpWYy79Rv
eug1L1b4kvRu7K8PHx6n7eaJgkIb+Ix5UWCwhUWR8DoZexYU2QShkE1xckGU4Cst90rtWIv16ByQ
YbMr5ZpFRPU2AtiYERtj0s65y6OwmVFfEp+Cxv/Q38viGE/QOMxPYCaxtuZ2/GfB4uRNVYNUp/r4
A+DK67SPDC8abmvY6P5ijIvhw9Rt3GVHU6gGeygGG637fu/0hQv9TS7CjQ3hfLN+0yxdMzwO2O4i
x8MpUl15dpUnWRnQkBxEnE3Izqrky/29t+/10bx6N4fZhhnwY+22pHUhhiVcUNo/Z54TvwNLTql0
Xo2/MryJZAEJn2UCbN5vmMNXnInDNeATM2nZM0gIjI4gS4Vx8LW2kj4Mbr10L0d4PdvlWCGBVKPO
yqIKXL+C7dKT2Ju9hn0Fq3pK3CtcpvT0q9CzVPqWqHWOTsxEBvqkEAy6KZnYJzV95ODoS6/Gog4V
RkO7XphwDkz2/MXyWy28ScW1ZDjGkAf9z6oNxRM5JB/g2xz2Q3CwOyyk1Fk3r0kh/njtwLwn+YoN
O6QTv6Y4gI54+60ijZWYlPrNR2VGN9qOS38aW7KPIfaM+iU/DXLYX/yykTBGazFAGuSKYR6Vp9Zs
XGJltsfsHeRnURlWFqU0JNraQFIaNAykd+wYlJ73iSfD8OX5byiIZq1gj4OlwOtQS7FOzSxwnyeA
GNW2M/nbOPDTzRRf422wmXvv/d5hZ1ZBTqR6xg85LXG2r5lri8bXO5gFCof+idJTb47JUkchK0yC
d6pmII8W9wKKhNXP8eEZd22DGLKQe8U0hmRV6zMfOQBKGt2DWCzPOLiyVVzDmFn9qRtvrzBbkvBz
658Dx1D/NVZoCG0w2Vhnh44vPxwUqaaME4MusvsB2cGxcn4qLjOju/aisy1ipCJhUwd1CXRqigVy
6Di88OP6QlZDpCdOci7gJDl5GlykEUgYiX4xQCdq2nr5R8uCwzC3IhkynShb1c6m8uSLdYE74uCs
ya3ONbiM9tLdJTRkhBfACxRoF6K9kgA17strqLP5hvnSt/G9v4UhRrtilR0U2QPznEVwVv42xzjs
xYZxsIG9gAvnHS8p7lheP5zjSjgPoVG1P1UK8nFcSvKXngkNoZ06QZhDi/AzuGRnQ65/RrTBkzJL
AlZ87K75hfpvCEy23soc9xLpkJjYRvSko8VgiHNgoN0ovyETBM0yXvv+z75FZ9p2kwKIAL9pArDa
onaK0e45eYhyhUUJdSsOFZd3whZ1yiLJLNWG/bmICKKJIzcytfM3H3cSMI/sPl3fPj/cHzvly/VU
wPYf2B2RGTrp6+aufbrOtcnwXiwzEAdg9mitHA4kcIQ7r58GqSCYPjOdVGHXYvReTpyAyFoBQCLe
SGHlRh2wY6gs5PnFCaWWUd+8pCvEovAh68ohOWDtlBDgmIyBjPBxfKhYKNz51nIWZztbGeZ6/i0e
VMgjyG7j/bj2SyNWbcEtHR/jCcxfdFsj1ZnmJvXHQP/xsynj6N7NDWcY7UdrPqQkALMdqAqEKOsn
UC/6lE8fh7DUmxQ3Ixl6HSmekurAZ0a+cIrs/9FiNXh35qT6Bs++y2eOGXNAKMLl1kKxEm3q62St
D51faEI9E8WhB9wE1kJk9rHAkGj9e6MJVpu5hX2dbdEkzEwnMZOISAvGKaAMWcGd2/mcBYpNcm6N
Slj/UT4Hx42mIltSf15R810a+3SQu6raL5FS+smlyIGnJ41MsweXmWy9Kp9mszV6255PkM6UlEj2
5qFItqxB+3E4qb71tjKFaf/qv/m85onUEVK8KPknWM74tGBMPqL0aK5xXQRidPURUFsv4Iu1ZnWs
kiedZvE0b/OMdJ5Bty+w1syoEPKKLyYZaa4KghoGJxAwAcnZj7hc61kdxa/vb+EIGEWVVZY901gy
ShVuBXlwkmQJyHvOYWQO0wjQptxQhhdUTeXAIZ/zUsteNEElTctorIK8bEF4dZUXYqK86wGzqczG
+JIwX8/OKQxJq3bdrpkYEu+1EWsw4+/MxJsetks3zhtXWSD+nDxL5OLebOfkxFrT1IcYc5CpQgbL
lypOCwhAz+biBZEo9OZXJsqu8Xxv45U1E9sU8BhT9SniEtwnUfzvULCTUvDR6bMM3ZmOCpBLcRWi
QjhndCg9xeIxeYNqblCiu/qjAj/G/QH3QuX8A+B71xHRfAxkoxsnr9RE+VYd1k0VlrAU3Q0hqkMm
pc4X6N07IksZRmeYiNSDXfcJ2npgRu5YzoIEzZhS9Aa6fvVXL24ARz0tiSOBPZDj/Uq+sBVFw64b
ux3t7a+xnMXzb2qcDGaABxLB0XJAtkIvRzUy+nKfRPj9JEpyMe/sm0cO0vTozyz76LJ4/IA/S4ug
ieiKQzZF4+s68riNzun99kbT4wstiDs38snx/MxDyMJLkUocE142t8LgCrnEj8StInVT4OKpaVuT
1t3dF4ZO5fwoRGHAUpVH9/ooBIrpVYZVN819Gwirk54o8EEQNxEBjvDpF3rR3GieLLCF78IXrP66
jl7XXmHbiPL8FVqSGtiy3vhUNQo7RbMkTTfyfp1QWtDKiUsFzJQp+9pS3R+a+lkxYxZRRAXUGfJX
gW6W99D+qZrdMsPgoOLbt303EDjeKb6m4foYaM8TlfZRuCGdYkuvh10f6mZBESr4ggcvMRv+aO0b
pV6mZ6SaNGVl+TOAY8NsfGO49JgZJr1FCKmBpy1nJ/bskiUgYtNj/1QR2ssUrbh8hC/nbF9B71ax
1MWAONHsqmZEpM6ipx9C5yvXrkwTpX9VSSulsSgXTGsGyW1Xq0PFtKTlaEE5iY4K4MlLp2Ucy5tK
yy35bhCBCtTg1DOikdQUVUD94naq12ADnuXTI8hti5zTJvb+uYh/6vqPHKQWfX3Womi107nLmmLv
k8CmtAySfkASeXuT9XXb/U6UY+6XWMGLO+9zgFuXoNqQv0mM41GZw4ucKeA0QIwu+C2aKmYSjtUj
DEbQuN0veJL3dylLcrCd+eZ/4VUeHjFxocGj65uW8B0v4zIuGwwipS2FEJi00Jd9lwOMMUJCI4aM
Qmpw3HWZaI8Sbos+Z5MNToPAh8I50u6nlROXUGK4fwok/T6YndTe/Qhfk0SGcgvIAwQMoftOSibw
IoBAOjXUNe5mfJkVPtr5e6ZD9GL4V/SjmRqIHeyj59VwGS9/Qir7vAZEhQggMnc6RevHIBAxLYXl
udWBPuv6WtYlqzgG1VbYt/UdBbfKlD89zAi2Cirr6hB8Ai1uG/MygHPsJunPM5ewHRZyXSU3Mgwz
4/saV7PT1CLqUn7bCAwWHeNMmiQWcniOTPsPKcLEITIrldwBBAYkFGwx+P0RUiIQg993tSWobolg
Z7mMk2Juy7WRRXGd2eCoyTByu7Wqclmf0LaIeS1SeXG6c0IqDQDhwv7ZJClX5U/TcEVpESN2g35h
coilfloNr073ztckVTEr6oMBR9DLdgga4v3dlQGfbt2D1KrB2IaESOgqc1yEEsi2SKyy2+vQ9eXq
UGrI2cj4gPEkMbJDWutL2keRWKU5fDBDZMGCZDs/V+PrNFB8UBaLNs0ttiGkHIDKXf3eaAbJmosZ
bji9bzuy4aN2dCpT/knbbYqwsZ7skQlgCyGbLLwclcPR0c9coGisVcfPSB8kFsCOXabQk3k7UtgH
IxkyivJxzPd/vTlnqf/RN57U5xqLSSwtHo9C5Xr9NoWtsEoG4eH55ENyWLqcE912tGSJQBN9Z1UQ
YDl/GnC7paI0B4c9AgGAIt4N0e0JytSPVSkyqfgJVRudmSZBBfZ/hW4z5PQ8mt/lbHktu5Fr3Cfk
ncFIp+tfnPXT4gei4uTY82ntr6HgYwjFSMCORThcKVZ3+Ee8Kxw78T3MvUzOGDd+uc+wyHJEe0Mv
NCjpaN/QYaRRffLeRVUjg5BXXg92PzV2j3IipVw2LLZeNsQ6OzApl++DUMZY8DgN13i6t0Vj3nvJ
d+wR5+95TCWGm0ZjNE5F80VgIj68p+IhitlMe8pjBum15D2oRr3L2/Xj0Z+3oW7vTk4VZuqcYtMQ
ABiR7es2LAl2j5zbfNopTOWi6PaeqGvxNulbbngEgbgxbWee6juVy9mnz8PiQmK2LPIk7jW/RIhL
VK0ikceq3jxGpF2DGx2dGPMiyuyvu3emTFd0a6G8Q0MNLk/2o4xM2bPNaOJWQyYXUpLk0l50ifUa
qoi19xLE4NzrQ6vAyralXBgeRv6d8+br6Yxco+AqH75sXyr7CweuLiso1Y4V/aJ7Y3XvGeZl615O
OGcrYGHB8p/6O1Fid18DlY0+HEI9zKLeoVcZvhUAghte8CdE3H6lZ4FMm7JQePxpJUvPh6xcOM1J
m3ivIEMEBqMcXQ0Czv4uSVslDLaLRfJqcJK8Js/RiuieyP2ROE9jUg0TavxGgHcUa6xYnzwTAU4h
X/ZKRIbbHJtWKWsUOEU8NaCCv4D96UzetlPZYGzgQuD+p/lO3IhhXY0el6WnP6HQ8UGz9QxsYekc
eQ289n1QM56WwFNE8Cinjgppkeklot10D7o/+UZvrNNFzZBGP2sP1chggsaHnYx89vz+3KKQp47g
UGqd5PyucWmGWeG9yfX268s11HZv0+zH9TD9k5a4fcV8CkaOrl1jgzBCBQroILsxCN8PYQ7GwXxi
RzAmnl83a+BC+isIpns/609VOWjbbbf/PiznLZclIBM7DKeO6l1W/pvOp3WhUQt0/tvBJWNgLqfz
RQnQ42Yzf1DcLRQuw/hNV1JH9L1HeMKgxGuCRZG89GXAxC+DN9sypRo+gxV4WSC0a3615Mcs5Lq1
z2YSPijn7LGzHC+cGBQggv2oR4OsNCkdKiYSbFCi6V4Fg3kiwBNVpAtwoCp6koWZeWXCvqoDJwbT
lhncbP2m2O+0x2XpF8Sbquw6DTrhmz3MUobfD5Z1sGpU5fMBJkSvRmA/9dO8o97aKds51LUu26mu
u/Hd2BGw0puYFrRs2lvCvAjwXJ5zTFEcpmRrRgmma4wWhOe2MN+5BYhv5DqEXmI/YHXlWt8dgaR4
myA07uhZEET8l/LBu8ZPDKMlfSlDq3i0MfhWgYb7v2l40WKXt36IBEY5I+IS68UXTzfu+d7rukZl
BVMugiwCrNBxSKjQzILfc8mHF2rup81jH0WLHF+S/kn9pYNsqHasd+FCAEP+7D1YRs+Tvq0tIEg3
/MSs4MxEqoOOSEhbBgi8Md43NBaJPrDmUUQPx63/RiRvRWlUcSfZ1/2m8A0A9JmEuIwP9S3/GLud
v7RKagHbk0AuNbSWpjIsXrvyifqcCpajcevxtcDtKd853E+pgmRVXDnG5VmgZi0BqcP2DaYUgiGc
0p5oRJq6bsRVlsXZyaZCDTc7pEsi06RyAwLqQBShDftVX/v0KHPcWAfEuYZLiCwYOPKIdaLSwYNo
d9rqEK99pj1Rfpql5T6icN4zBrFCtW9g1Nko6e3i3Z4nB8YNn4S1wL6TCSeKu44QKV4qL14TZGma
Qq67hdCb0Y+4v8l6T9vVzb80RmT1NbofhNeqyfSzEB7Sb9BRnsa1bsnWFuK5duTHfnL2STgj2MbK
6JqtBME1iwEt+LZxoCxC7PECEQjDd/zLi2zjfHdjlFxSHS2PNa/WUSm1hAhejG2JIwjH4An9ZTD1
DIKPvxDG48uWocJKvOjzmPsCSJt8xk9IDzVc5XWyi3WzDJA0lBJr7vltJFXiOabMv1LXZBUve5oU
1aukA+Cj1oUIzsnIVcoRGJgUeQtqJN49i2tGbbsXmqNEHJ2BIUl+XNnOMmRnIBK+1DBzTOSL/ZQh
2oppuZdm0HF9VMH6KXvyJfNkUIChBGWYtv3JRbTiAB5s3PAxPoSCGRnzyj89iHZw9TQ5/0T0xiUA
0m8NRoPG60irIHJcy79hl3y13E1RPjzhTwUuDh2iQ1Me/3UFKb3XIhXXznSZ/ryhlCJHqMV/fePV
OD4jydv90QaMrB6/Kpy0KtEdBh1/tBX2Ndvt8iNQra8+A4Nu5Svv0iKKTfGeXvis9e8UQrKUwjkw
wRTYMRPxAZfD2lfqovTy1ZVEj66mE7DJHBp7eyRk+jv0qh3Hhn6YFj06MfbTai8qhLRyhI3ojjKA
LXSCUyIN5dukfuc1/1R9pdCt65uMepUlJEcGnFUjLMeT7myLcKdOenrhGW24KB0M+Of+oArR3HB6
55pnXH5CdonvPUnhTyFYSu/44NTW/gENaBjFhedJmymRfQkHgsGhfvEPh7kbMp4Dgk/NSbjfB+bS
GmtQeUQJgPOiZ0Pj6CbHhZjJixVqGp+QOhhT3GcZIgs58Bi3hVx902CiC9XmTB3d9d9XQJcljN++
k0Otwv+pYX1qRGe+ZGVmfAyF46uFuNwEJppwFMOTsn4SynQLyD3FNlBcoUFCq4s6dK/z/waxcZxv
LQbGtqaRa/68XsELCkRAvIjqPiaVfhugMaHOFkrT2TBoDFLG53WTUJj/wuX6H4+FrHpbcItRmkR5
8xG7pbnt9Zc/GYg8uY35key/BhTfo6FatLcv5dbDXvCBTSY6gqmSF5pQ7ZkxOpsows2lLA/wRkFZ
0q+4I2vmWRfjjyrNK6b9e3Os8uH/0pCnxirQWLBCd91S+9E6yTmVqlik1GLqU3TheFWwIKl0ZmP2
cFafGNL6V9nykOOGmA5phDEjd4nK/UxJhmk4GsOvVtqQmg+KGiT57kvoi9JjGUwn//kbWdz6cWAx
kpUEadtophJOF0WcTuzHDw3fSVJ7YCrWcrhzBzSLFCdpiE6raHUn9zsQ1gMal7XUVHbxdQbVu2CU
247R1RqJIBTUj858fUOTkMDh2lPJ4+90pIcXCzHYgy6U2xj6v5OZSQWesR1iVZ0Ie/ayAKG9/zWT
wC6k5JeyKfMeizRkNKRKRwS5pXp1liRidUOZXHHeQhGHoc3/DVZ3idYHxmTZ++uv4boOUJa3L/8T
KZeUGVK+tK9borq9e02jtix34wUN4u2F8WhK6TWy5ocv5c9+kBcgpqe5sCN0gbAkME8b5JLrQyED
NGHZPcolCPOVgI3pkrl1/1kprU9HPJ43CcHR/Shg4Doi42S4l7OsYoZRmgESgPexRzmrAEBYFZp9
2q2bjhMv0KbTM8PSpa6mAgWLeRuZJ+0FJtdvpUA/vMZiRduqJxJ4dLz7SzVKwhnQKuotaWsMY3TQ
rhguulfvn88MbiTp94emFubbWedZdLCeq7kRUdmL3rxYLn1zWqZUwcOrtZRqTKalPvXbDJAC1e4A
4uPVnJGw23AOpflmbfkY1x0nyEGKGIpxveclmYuGqVEbBpZ1vU8uO4m6T6vKwj2StaMKBTdB1HqQ
tnOzb5RtMdQ/WwOR85fKOcC1DgOpM8ZlfP32lCqDrM6dt13Trv41Z2x4VEpak8IqUSrYFF65ONud
Zed1/OI8Rob+p+yIe677VnbZUixhnx+PXCi5n2bqdsTs1ZgcR7Us4Evn7+HkS24MOVvlNc7lTsv7
RbArunBSiDKS1+5Ayp5cGq1qorf0qYILAkhPI7/seX/OgCcon/7/dKVjZjSxoioJF41S9s5c2/ZM
3D098vix+EYvGnxzRGHIizL6MVVnXiAbvQzdQR4WULu5TEO7jSXn1OF+K+NA5FrwRUd3TRec/jtc
J4veHdYCJa6DT4D++b0qT0pxen6uSHR2JwPUqpzmw6+M1+Zv2IyY6jSzWCCb5HZdObXQOAXRTaWo
Qx2Cn1U0wfrWklI9t9FcMJA3olKdgJfHbiNb4FEi8KZAsdsEkuW8UPthCd/1Jgd5suEXk1esLcM5
Ud6eFXRhY9GwUGcX5Vj3E4dVHA82tb9dxTuQM24QrLKF8rDnJzGP7E0s0Lmkhx1KAOKV+BWlR3i/
Gh85uU0idRk7gjHOTmi8sDDNTMwR3WJJQt2LniGcS59f+Ej3Ko5AMQaJZOlFxIUwsxXcpTjKX9c7
tNd9pd757EZQ3l5H4mxZj3Zf/uAQSK9NqPDhV6aQ6rLDSAaHvqiX44ufecR52U+gR5LFo233ji2F
ZfCfg9CrE2xFTQa99Ytumne91JWrSL9qMyGKnTr5dTWrjoEqkEqDNGH5d2+iyNce/qZkeTSfVBKH
oBWwpjkFB4z6HM+dfowE7RJ3zlE81bJ9R0gdZIv2XhQGGIw4cXufCXPNM3ips20Dp2s+UwRtluEU
5rjOxFKHHO2gJxQS9VneF8xN0q0ZDtImwpqsNpLyRAJDlBgU19t/bKXWecJjfArzztdslBPQgA00
xsA4HnXVLKVWeKeh6B5pTO1LrjtfuOpb2YiGnBBMlqq0LMKcNJTk/UQNaWCxFJTbw8nfruHVvBEa
wyMQKWfcakv16tqJwiQ7OVkCIbMO9ydXnG4UdsorREX40EH4sbJUOAgM2QhYOkwWxHQa+BGuejG7
f655+sSRgenYbr6wVbC72GCp5QyUFZ6YBMy6Xl15GTeY0r6O8hmbJmY9rll8Vi3acvGlTSLAbVsK
GqkKHF5VadG9Jkds4dGxpRHfJjyirxACpy045Ma6f5htpgLyetY7mpW2fPgGWZ4K4D2AHuQ+OVIH
U5SCqvCvdOxk3iJPPiusyX7KGNj5G62ipX2OyRnAJIjTSHMtIrXSsw61Fo1NeC57dMG8BezCo+N5
6x7B8qjeHjW26xdhJd+JmQmN/DMQGakzXcsLBMbFxLVfYhzp02jVag/SuPLIW1nf5u3zZl7NoX2i
YEkfl/PgcwJe9mwZ1XWwHU1lmwRKkjeiyEafchlH05zmOcxv+DaMJdTdEHjCwwcIO8Qi8Tb/1lTw
DUQBYB+SrVqDHIXZk24K44Zc0/Ty8YCZeVqx/qgT0lmTqGbukfg85EVSvupvJykJFV7BLIjS+KV2
LOwQRbhN7hNs1ZnjFBbldA92tSU8p5zCqEoBd7d92YtT6pGCOCUVNUnGoRsXRKmu8Tl8ph2lQK3q
EBrZcj3+loUkbX/P4uAVgbwfZA+rViYcSByVEUVJRRypL2yNVqaZT2TXeM1WWXH/zlrOjTs7xvLa
zzME83ACZFsPA9O+Y7GEsQahRlpoHmT0qPSunkT6B9i9psjGVX2/hDNE3zxRW8pNvXoLwq5U47KZ
TU63L6WGe4CtDPFFPXZEHT+Rpoa/moRiEAI8AvS4HtwYUOFVZdOp6ibD195UirjNFUpNSVd5g1OX
2ZrTzp05ezLbYM22cb8xWJHDOfbRyaj2x7Y0+bBCtBRqf91eAb4aN/wHrTgbae2FZnxyKnDHc9Nd
bdqzMXwo/ND8gMzi9IAY4J9ubSMmVxBHk+9hBr93sMIQgAuAoDB2NpsX7rYZkf8fj1xcWug0yo1w
TjV4NEPKMTUbO9XJp2yjOuZUPc36HkS2aM/IStrKXou/qXVu5wtnzBF6R0J1+ptucWGFRt15H7hK
t089+hGheAv6tz9L2YGMVOkJjWDrYgKjaoz1C1sulvLyyyCbQts/gNQDZcX1ONucorhRxs1t1NjF
ox4PzUMJ9e5I856lrfdTWIeYtM6Z0SeMAvPZIzlIaQvGL8UtlGyGYC/dGzG1qFhJAD+FOr0wRUln
94Uj9JTINsa0iUqXDMYRtShIdNRNUCAjSTN2B8Gzsz+hgnTzQUDVrVzVcjVwG1xypQ4IHq8TI170
9eDgst91ZMmwQk5OA64CYOYUG6AibBDYIicy2HlZJdwpmjysPM2m5V4XVViVHYbR1xwp6ASI8+hZ
0QZOj967euUdQrwdqScX+bMr5a9D8ptFc7h6eiMVLeT+K3PmMNU9NngVLUgTdeHWcbWZxV7FWrJt
9TeM+Viypnbxdng2GoVGpZtRKt3inDnUgvVvV5wMnhZyVIo/lxnDbvitrccVP2eOt0HpXLuj3NY8
TbmAAozjREQn6bRlkA4oJbUL3DRgi5Fw2B7byB2+1/3IgBdk8/s5HTjD96DRxJP5rI0XzZKE8yEG
lHd3VKZv8rKF6fIvH0fcMtuR3Jf+skMHvSk23aMAGhW5he+XWLqYTW3ggVCClMDuqq1w/p6QdRAk
ah1sf2Npcik3BxS5V7iWULOoxX8hbfRYJU2A03hgVBdnR4qRnbMCnkoUi38kxFw8e4XTtLpIhT8M
MGHw2Tjql9I3kbgUxWYNZ8SsK8g6Xp3mj+pBap6T5oFkDuCtMU7IZVa5OcyAmpdwjhQtzKwFnJ+E
/NlvlY24jR3KJ3TBgCAxGiLcPrcZ1N59iL0dwxz8AVuLLCjRihUSIR8XvDAhJxizwJqFznWa+CTc
Q6Jp6TwCRBLD9fvlxVhuy6fDalS7CIFiUytVzcHHNxbXAuiDj9Dp/+Zb+9I9IfTzPlfDjNUSK/3u
+TwuLHIYpuxy72MvlyuVX9Xxigfu8nWqlFzQkohSFgWnaTC/eUWwCWCK3n218xqQY759Gq18sDM+
04GuOhOWKyPMmoGjZmgE+W0FdQM2xXmyrHg0tIz3R+1Ued5Hvj6IPFggoJ9IGNvg6LRtT6mLVKJM
UflVghj0GabLe668Xow4oWjtH6sioBB73I6PX9IVSCQg1EdLZ7WvHLqiBw0Uw8mxYFR19BbWI4Ks
F8CFkjXA4yIp72EscETwoi6il9UrpowQNGByKy7HvEYcZtO2R6iihzCdY8Zy/doxo80ak/wRRuMN
8r8SpOwicERlW8c5mb3Dzw4cTiHt932MItv8cjxEIY+v3zZ41QA9Rm0hbS5on0V5w5Wdg8MWU4cT
qjZpvM/MPLIYCpNstUOc0KFLLsef90DQvGvOhBnBsrUFxeST6WX7PTQl0ava+FW4jtB9bDUek1fH
eqpvM0afcEaXJNAVudOHYJnUmiEZxSLb2LJ1h9mfopJaASihl7TIdZrb2xROeK1G/F54BJev91kq
CtfTpWw8HL3Z/vsKpvZPkyixObtJlexxf4h3tmbw2vrIa9PZJyrBZczhtYdsabdiyeh8RDd3vzVO
rfLQQ8HbY9HiTFv2umzbGTS+BiuucRrr9oZcCxwmUIt42bo9F9qFHbJEEni8n/B4C43RJonP+y29
Mp9zeGsXCEQizsx9ohsB9b2PCGkImJOxpMw4OpAB2M7q5T8Gb3vxBqxViD0aJUa77woqqgWH1DWX
KnOBaxYAT3FcZEvhCGLo5DRGLPfOzGmYb6ysLaKyqMc128Xhg/bZMp5UoRB6+dccZxgbKPfJ4n0h
bGYjO4GRZnNOwb9Hic5SjeaYOWhvtORjbMGwCEWkhOUKgVVUUEw8ac0eNWbVPm0V5K5MJa8cXTSA
jkoWlFhMUB8DzQ0pjyjdkfxAFb03n7Uw1qbLcd+N/OQojrMNi4dzTaO2MQpC0HBosMVfJG13igBw
z88R0myu6JJSUPnXdw+iME0eeM7E2DtOeDBNpJPdlgsPguGxXdjqsOLPHdBtKkondhiEN7IA6IiC
xdpA5Ub5wM5WmgODl1qEnAFFUUSfE3uQdPL9kahWgwKxt0uns36J7FJT+mVklN4r6kEOLF4FHASA
koNhQYsv0NRcifLEO4DFHpZ0l8w1wLmCil7ZrVPAySuEn7ejKHUB3+F5L1+SBiWf8+x2vu7r0bpq
xugN7DOO8+vG/JZdUCcueJbtPgddj7nJB4A56Ie/xsbatkLIzVJ7UZjzBULtTBTLhaNEpHDyKoof
at+hCOs9aGQkVpHHM0vmTFZZBJkydoSR+zVWe0C0YgfERKXgHpN+4ZiOnA3TOCWA1WrIHd7Sx7SJ
jXfKCcdYnMQOR5lFUi0sjbMbwUK7Db1ilgzCIJmSv/AoNQYYZpxbTNl5bAJBOOpmHxYiNI4U56MW
cs4f+E+BAdS9GnRmfMltWLGp326+DznIEq1qOPVY769JkpRt/Ew8czxP0bKLi3IoxpLyCl+EpcCo
Axtv59PX1ljQsx8Pu/66K+h1zcT4WKo1qnJ/BvKUubdlsJ9alqBH4V+oiGQ0K9KGEYvSRTV0YWNo
ZQkOO/IOsZwVa5++r74GYTnKUCa4m02TFXFGntkn/Ld0fiLiuu6K2oMg0gUU//hP942s+oAVMwL+
yXE7iO0CDP6KLqFqezM8b+JMCJExa+sQY5MjGEnoDvE1QXVHpdOaMD0gFVcLzPMfZkx013xloGvC
43VJrD/F0MoEh5mPV8tBp13XHH/kWxmHptVvzdQrdEl75Dh0KduEsDp86EK36ZAEhWvRRfy9YXq5
abR7P9/aXK6gMWRQq+J9rUqXSRV/BHQqmyiL3y0oIAPE3/oARQsvnLXJYp0aCM/Wf4pV/jA9RRfZ
z5oo//5zFedKxJjalhchz56lbR3B96U/zks3iQy+Fw50hTT/Qagim2yFLt9oIRlCcf/vuLtXLECI
rb2H3a45rCDgeriWlifYZTrROyw1XHkk0lvUg6IaUYRV4BTwz9DefdJ9DP+RXMwbc3NexInX2I3c
fjsPb2vt4kBo7S1jwhqb/i99gDcqs0pf5N1cQ6T/xOuMHwmk5gbntBwfYfFz5A3WFoY9BME/4bf+
aBCClB7mQPo1jDBonflJQanHrSxHq0zc8wLi8qQz4Rb4mcS2dYb2PY3Ed3CFMCqCqpkpkWgaciHa
eEqgiJ2ld4k3bN6w3XhWe3VYkwY3mZ5wyFJnCfuXsVpGa+hhWq5efqMmyY4qA93bRdhwiq9FQju8
jWQrD040wRvwb1PZsCZEP1ctx+I98UJN/ovYqLNGgZ7c02eqaBS/ZU4WWiyG1M2cmcP2pDhbryUd
BZZrb1UYZQWQej7JtTWW9Pt19Oq2uf2k1Z/NlyotH9g7mHQZnWLChxZ1blV67GUpAI2KXRi3VGb4
R27ABQ/5KPTFZLweWEcAjEER/4wmlRCD+6y83LxfV9RyeUM0+/xRbZWTOroB75fpBMLxE0yIlo04
VeTCjxctMWxMUxhD4TMF9qMq9NQ+zPdbfb3cxSTqOiqPVd5roHoyWadA+uL78mNb+EmJWhXVt0jU
muzJPvZgVBgAipnG7Wa2xEi342dvZxPT5umZm2FNkJwvuzlUgp/Pet3iobLQKq1mQZbEyo3GMeZW
kxK9xTtbif/SJ1tH1FsfmPR3OPVB49NOWJSWeNB0wAllfpo7hfT4PpPYouxZ3iM2MTae8SqZY8yh
9tQjB2mwbzKdlb2NGr+oPV7LwYFK6Eh6sslUERYBe7uJp4zL4V4Xyxs12BqRajDlMo7zkdeV3RS7
uKNqONvjDd2ixKhsvg+OkW3HYor3kPVnbOsJX7KGyLbuKVDl3gtw4zZ1Z6qxp2wX6hUWTcO0V206
NVd1Sjqq/PQWes+ICZi8NTv/4Ky/ofdKRfABFO8BbvcSnfLq1o/Ryoe5za5rTA4tFO2xnP/3iTSg
Np7/WvDwdtiCXfFjX/vPWlO3GJnh0q//mGQg4fD0ubXztpuCdsCnp76yyb0up5Pbn3l4+Co3HWll
cBJKTK41XzFmZTu6fOGKOuF3tJoLHV7DSZ15EdRbRdzRdNRwP/9jVpycBTAC9zgWkcW1rN+u0/4I
WdkGh+vnmCnF3c0hg2Qp0hVOR/n5t9cDwyhLUUsweCZ28FAJT0/T3ekKvIwWXuystAGJuqr1zdcH
65fvODHaOLqC1l90WdqEEy17jKPYbLfrP89vYeRh2cjgsZRq7dQ6tUiO0tM0jlVtPnERPcBdqAEU
5y82/bxnoiKp7b/6w0wRhGyBuTF2ExFKvXYsV8mimsRj1bdHpTeazigKDgQOkUcLDAXBBQhmtG4W
swpNjFdYZ56wP7pnB4eZnzd6nN4BiOJeYgzTZ8za4lG/FoOm5Yw1o8tP4H35nhWhNeRiRlYuz9vE
yTdk70HawgHGZYBPKxfpXZrCwMp2qa+EhmjyxO8cuiIwQpd6jxEjNNwmzTWvSCRxeEnCxG9hNTWd
CUvUv5X5EdgyRhAf4Dc1I2hy/7dI8hlVGAi+orDQqyfLVWF2qmlgLfn93R/P7G4XkI2fBz0RKnQV
IeNtNkpa2JIEoySwqstSL1wVjXTLyottfuGv2rLi76QmFy3ORYxXI6Vn3i1vGpm9tKrnMzTScoDp
WSsJsBghGmfs6Px/l3KLzO+Ab7ImB61tyqrWoUAr75l4DsOAuI2oE03TFiePtVnzV/nZFOq1tR0x
XaZLRz8UEF2loPF2fzQ+K7f2d1t11cZmowdZoe5frC2P/pJnagvE2PlReRsKYHdSQog/Da880jQw
CRz7gpDBfxvBtGnYQVDuBTyRPIm8+j9WNE2giYznxTu6PJHtspM2KiinkTdEhALtvUGvLuhrXkOs
viuE2DxYGtt0gQltklgV5956vMJgOQ1PJFe8UfXrDhRvek0LFlE4b3B5jR7faOensJai3trWA4En
ChVe2j3S5GkduG3/pliwauaJgtiKN23w+v0rRSbzaVug9v11gi18oE49AcFUv4ZTouSIyi0sVecs
NlouFKUkbCFNvT7pOtJ3/7+qh02Obiz7kUyOEl8EsNS3PADefJEUgZ5lSDLp3W7vFgz4wBgJXaX+
wrlep6iNTGubjxOIy8T53zzPLkb2KzdfQUynpRuLOarlyQ8SJuf0AOCONjSWpcoJib7AzmsZUfxb
VYIJ3nmffkrC6FfGZDMkfMzzGy+yroexFoByZFSLwAmq17/w+vRJJMnl101HHuokjRGTXyk39qOd
YjK+JphVvaoJ0+fy4jVzEGen1tNbjUI4F560y+g5epepQoUSGOOPwnzJmXzox2pfxVKzz5V0m3hQ
F0bo43ybxTIzmXk/GkRjOsnHtS+jhFg5AlehTVnMT8o+ct+J0eDTWMEvROp/KoJttOHgbrtJxzkY
hhrMMIEISUpfQn4Rzg0drSu2G68CgiQWYo/quDsrBKUGQgMOago8QAzc60HLH9JDZ8rBshZGKlt0
q3t0RjRcUB30Zsqxteqqi7I0x8BVi85cTY3IfRMLb3BQI2MF7SWmsCY1AHhmJkvr5+GfaV/uvHZN
zRTNytvCcd+PYJ8qx4uyk3bL5Yg/wTy0rwfs63GyXj0Z/iWAwyqWqeeG2Gg0d7KZZSsVytfqthBK
hmd3YTRvYW07kcWzLTArOQVCDAj+d4LF26gNx5z04NJYbc3s3xsPnlIwnNCfD2nXapVgeFmkLfZY
CXunWXXtVXkhXz2ZEzyjcK8W0a3ZqF4j/7f3Z4o9UMMndocMv08c6MAdLWixP6ryko3JIlmfQMdc
JpDtP3LrMQUUVbCh+S+zfB4p/MGvEb7vY+X+pDW8Bqm/GMD4cM4McOqM102e1Ph5p+7hxthB1ROJ
66k12GjVTwHOTGrlMX2mTPjKandSqb6fXz0SSLgUA1iU/9jKT4osLy+NI8qQvSbmhXVMlUU3hLs6
d0uiOx7rDGdk7GPsTQca8062eLpX7G+6ZrDVCSJrFtatnMEbIpOjB3Dz01m8igK5RBUrYgcrn6D2
GpqRE3sKAgZ+cN35biunOyqjQQqMK59NIYnjQYRpsbJGzG890LUG69MoBpYYLAt+02m23sU8pzYX
FKgkEJE2hkwTBGCYMGFmb7sAWoErmzgC65iADAEiy/IOW/x8bIzyc+1VPgQTsYNvuWVEBpbgJGec
viXwBlc5mw//9wxWxE/wLSeBvTzwpGYZAKcKGkqiJGmYCAV9ubdn1QnBVMGYZ+VAHVh0eUCAcrDJ
lsMKB+4MH5gpk/HY2NKAKPCULnWgx7IhYVE7DFOT5x/L5rH5SrvgFQc/TWj8QZbscAYQOsAiv0s/
Dhn3EjJho4cMU6tbxLvPijLiWMgR6kMEHRsylmzqSyqsg57Ht01HQInIwoc9VtSHScVQOUcOcDP3
qz8wH5b1EuWkHlKq57lHKtNVwxg/37qrwuDbsKa7B5/ZAT7va176ASQyOaBVaSKUKt7IP9b9QO8D
gJ+AwxhMKx9+4mK31ltIN5hXgIIy5TBpAUnBeJHUIG73AO5+iFutuXLWYj1jBODkarnrKC+u0Rg3
XzBgdQrr0WxNC0Poy5A8G+oZe/nRYUEfkdPs5DlJulE0xjvbeeGxrl/AAZLVVO8Q/8eKckKXTQJ/
+Bq09vPLUT6PueovIAwHCqaH38tXAYUpA6y4c8wUPnM7zi5gDFl57h2MAYcHS6wb/oEycyQcEKSR
6Nc5jkwGCKZ3+4h5p3gkbhrq30+NE4q6IqEDdTODrLoqDsaWc2h98wYNDSU8jJlEWBZpRmKhp7O7
iPBxydmsltiZOuuP1Jz6hNRFIScNc+exwN+GG1Qs7zNizcXJwFJdV4j2DMynD1SmZ8r/YCT7Jq/F
hfDD7j0WgdH7zE/mG1Y8KvtlJm3X6R3fdH1FpOFx9EAXFytjlbYqegntxNK3TjD4rC2+m5Y3GeVr
W+mweJUunbuj/EdVNe0ycohXJCY9vSQNW0h/mYFOHlPNKnB0YzWG/7Te5YCqgv4J34gx3zzvbLzv
g/QoCYELpSM+FQBmDlhoBS3LHxKh4mwA/Z5/tfivuWbUxyyhgEGoixgMGn3Pj27fdxb6qnF9H41n
2rru69sbYakv208NBozfObzxESxGJJTglEQOxnYW3OF81rnpxA9rcg5lAA4wfgUAAyZqutiQFrja
txeB9pg2E7P4vxxhB9xJUW5YK4VbYfugx/A7rt/Ee+VV3qbPtb+VcQ5y8Y9qI7Hg+8Xz8E+prILn
JZ2VmQWz0Xc1AjLRUsaC9/wdIGY1YJoZifo1JDAA3xRVZ9/DWEkz+5rd4TiMf2Ca7BxKVBm3fgGG
tMM3hMU9V2XK+i5TMrsv1aHJwDw0q2DXUiETjxCNFvXNV1RAGZr7BR1g+F6/vj2rIcXlIMy+jJg6
dECd0kTM560RyuSQjU8spcbPwl5wGfbpoNRxFVIcXiBUbF6QWk3zDZfKayutKg7GKQ1/MCJh4D3Y
LUE9nhw4YXT3lsnbm9ISOqqY30C1+HaJs2Gfx3t56QQbscfQ2CvWblMvUsXgY71V295fhjVjYNxb
EZdRPMnFD3iab4qJYuBGzEtBUOXHeudW1R1WBApsun9LeZLXzri9CqU6SgwVYOBEM2cKycz3XO8u
0e1viSV2pdg3ihHBxtJoTB1+6Pj9mKOCfJi81fYPrIQ398Mnommf0R/OOOMu8aY28y8/oloBzH3Z
NPbx1Qm+4t20WzQItePMGNeXIQs33xe9K28++KD7/UyuBqnRM3rV64wCUU956q1dSrrUBLRk6i+w
LoE6V5JaLuxT7SAogemhuB6BDeMdeAxJIbKiVtrfsUHgYSmQZkDJP2cFpSIBpXwF6D+Y14J5Bsqk
GOn2mfQzT7ZBfv3eeIUDiro2sWL3AP67t+hAW60t7c192C4s1Q0XV72p4hR3yE/t3kjyTS5qeS/O
yl0YiEXe6n3aZv+nDCKU+r3oJ3AgRTPvCoIDGfh+AskSozghzGToiatoxXPVyuvfDM0QDJBbuBgf
43EG/BFAiBARjmgmvOBrL+1J8J4qTHRq9D2ha4ZkkC+3/G+M0axoSrw3IR0fIkDQ6owkXOYr8pd7
KRdOwTFIP1GBEZoG8Wfhw744RV/MU5H6uDnjlZeMXO7ZLswRcL+RR580whVyz+pMBQcfXJGOOrBI
3Zo0CXBVdUX6KfngiU04N1HH077FHf9IZr/M5aLzFIf4qPHAlWhFMWY/9Q3bB9updebRW8yExwMi
UrCu9q9PYEmUhuS3dbX8t+KjbJ2RqMyPuwwxTwwvnjYXFjVdCmQ5KKlURO8ibEj/kOQrhdT351li
eKBxJZ3zOsVVYYgWAqmODJyunafT3ZhGG5HuvEwMu7WvwsFz0frz2QyYXNv7IruwNHjDBQA71Gel
xaP5d9GEdTh884BMgpBfbBgueDbo0G2mzcFBniKFwfkqaikfWtU8OoirOKpfH1/N8Qg4CMiOLmOu
99U8PCXrjUdpGM5uB0hdxOPTN/Ewq0NA0yFs9I7GZdkIX6QCe0ylAkSpwjbLglxQZcUcap8w0MLw
1qs8ARzLdqF9056/wyStCd1pIEhseVDkpxZhw7RAv68dKR3qclgewUbeEmSHNSwE9FR6S8Msajqz
kexFJEQLOWe9C+ANnyovx3yC9Cj4L1jx1lRy5ldcNEjVeUHm/nfEb8G162IeGqBniRcRRVYNqGXg
NJCeUDZ8ajUwB0cdiejsu459Z4WxVSEWrB1mJo4To+ZmgwW8s+uzv63pxx2bBHBzJNZ34ZtQwszE
7eP8x7PHeGUDp1CANfXiM/tQboKdE6ufVavVctt+BKjjRGBiRH7ocK0ACfIOS4ZgUIDd7biAFWJd
TpBK1NG0E11ALXIhFS0woLIy83G1g4YiewFaeRuq3q3pMUdCiflCC4CJMi3NVlNmfkf7T6ERzi/p
iM6PDPmfejWcESqVBURJSpbtKXMCMXDUV4PJM80NBO0H7HmGulbsSa9t+L4uxaWzQcFDcgitI+bI
Ipro1tTqCSzDoSDo+/nmMx2V0ZVwUpgc3arOdlobD95pG9DrmxpLj2X+xVrVFpc08yZJWas7uLfd
0dJIXuI6e+7vgRQ6ZJHLb8dBqmONYPQonfjLfmLQfXmR1WIIitJI5gPVyM3xfCFKpFL3+yGQ0Xl6
9AYourCVNcJUIZavZ989jSAh2nK39298hMemHvSMlQ5wgy97KrTDgtFdb3/3HyBW2hWoc9h0tsJA
piLt+HmAPM8jNOMFG5t7FilpZS9ES471n/nr0S1MIamm7nGaQKewPEJqR1SFVWg1a8E9S3qR7Enc
OmjvEqYE2xGHPIrDF387npxm2UNgbOXr1o9i0TFTasECr8vnBKDnLiir+D1hxrkkLaCOoe48a2wi
/AeX59j9024AQGCSGyRQ478mZvGnWc3YKrwk+SSHAZOTScIS9qq2OJ38A1vWPzwQ2HDJmTfXrSGf
QjLl2Dn6QnWKzcPXHjgFfc0MUXVGP7vjX0nhLfDjiaMhKCJczlZaD/yyvUxV29I082Dk3MseXZWD
Hl2aJUw2/NCOLp376M94VFUr31zKbsRYqcQyctfFgBDKn7tTry0DG2QzhjPTN6d73eY/aizwwsIO
MPXpUfI9b1wFSwlsgnMz8EsgXqK2+KpwKEW4Qs3vLad+dAQsBJ+Ig88bCqHERPuhvQUKEex3da+H
aBbL3Zx69JDUg/GD+gwIBRkPusyYTS1XzkuvXbQ4fvjw05vSS5bxlylkxfSK3/ntc6TLHDR59l68
60LPdxiZnb15wTF/rtlo67mPE2UsOOX+AeiOZqpixbk+QKFkuASai6cq1irdyolVqpeleFA1Gk51
srn9CDm2gdIqG9CxD5vtszqxhWkMKZCQrFe0XFbr7YW+LEuYDjLBBHJIUH85zSv+yyAm56/DJrEU
gpA2VYVc94Brt4AmzSaWojYa1AUyaQBrkexrnHibb7FFuC7VIcJdUJeO05v6+8vawLARTAwjNktI
ZrVgwwUBP8qyOzY25utZqMTsVwUaQWEhVLtrRh0Nmyxl9Qua9mG8Sbw+9AKk7gU61Eyzshe7yB7c
Xk2FpVbVx0umqw/ng/7FgK1gn3WGUcFmzkBX2Okf4jEfu3ok6zSyCntPCeqfYEFAM0bGHUHyGQ9U
wjaKJt7xSZX5T9bkR3bJBnsKXS2vwDfrGwAqi4K14tW7ERcKY1rlwZhT5qAVigJNA/w7U1v8xgHZ
uSBIw+GeBunmLQ2xdBcibmi0Ctq7EWIEvW0VjL1r75NM8LrhZEPNTx25BlEIZLB7PH8uG4B9YvwX
mlfxVGmQrEPdqWSaGuNEonf2kVxFuSbN4suQLyR7os1nDPZoyahQTSH+k9vlJ8VGjzsxWcxbzUt/
0wrP1+M8lNAmCsgftpyd2SiO0Fh0NRAY8f1j8x00LUrEXA9muTnKjA8z/W+BmlgKWVEBYsUlLSne
Ej9cb/efU9P9nfybHetofYt1CR7LIk7tn8JmgQAgOQJB3FHc6n6r+Xaf5ofbySNm6Lj9vdKgybsm
arPr7O+DKxMrVP6YyTA0Lf83aEo1PhjhyD4tF260V/i6Y33hZ1IjTxzkYoQO4qZp5lhLB6V/t028
MIBUSVbBL4d9K7xFcLWULVmku+n4vDUmv38YKq2bJMSWwlwg63icu0NeksAfJYrdz2DwcSmwlHoM
/rwtcCPzr4SYduXy3GLvkmEA6sbP2XRASJRCZuT458fa6bnr0XnXVsxFipv5mGCmoMDlHx1YFA0x
HbEeAPvySPLzsbudMTRMF+3HgIa9x5TLJLAGpFrTTsCAlIpKjm05p73//wjwykSjcWbdYWy+h795
hm/rBtQChlpGR5RA1qa30vRdQ8AM1lVhJF8QNX6eHPHckENcaKPRYxapISC0owNqSePSpLwBtduu
BSKaQmy0EV96bcSUAXrJZY5nE+jenAtFblCT4N/WfVlRop+XaXlXDUUWygAgKr3toN747rKsx5La
nR+qfS43IbeZe9hW4nC/L16PzBhAdXMf3pRSrEbZvUSzwhrefYVzWN1zcFaeOvg1x0rQtuUnBiVP
QVd/F5PLYKc3347dJ88Q8fY5Dy838gHegx4CyMfWvgvODgBxWhv/LPEB3PyDTWkEjuiJrH7LyAPB
4bRYbCD05vkwBVOif+o7FYd8CrasxZd2nDbZVtQjeNZhqgNdQtDSPnFV4bd+NWPi1/CCSY+F1FzN
4ZZpX/aftTI20aIz4DttOmltwJ2Ccv0JmrQ/hHzOvCCk3T84gSFPPxMJ/iFK7XPzwWd7xyQDpYSR
y6WQiumQFdAXdI4LvMTJczocNCNx/0z8VzJESkFVHR9bzqorOqYb4JYBa3bdBPn2Tg+pdJGAZvTC
XiNwGbz+usXSk4JeZM3ggDHuwwhcN+3j12A4Q8RuzKX0j1VlMN4d07/KDo5SvmLtYtBcCT1iNJhj
LfyfAbE2F95WxdX3yTYomK0t+2jcYzzp/dY4CHbqxhNO9rapn/T8Q5pCLW+ZD8ULTbCZ9UfGJzxf
S3NFdUwfxtyM1OP0wY/HjFPqiA+wzqNhtFYk3esOO2wty2PNUn1mUaawgbjzm67Pdc9xHIeqIdvW
e7589aS85T0LvSE54P5HXrsWqRLYhIwl8M9ck7wCT56y7o+N3KoOQweJ3XLP2LH0bNu7fP/5XDjx
SWZnFovzKoaH8BsBKIdvmTQ5sxdocPuAWEx9dFfG1Nguqqq3/O/gSY1tT0a5iY1rd9OwMNBUTLZH
y8u5PAJcLjagxFsCRlAVMcqOmkAicacC8mZnGwkN4tsejz88/LalH3uFBj6fUncq4lD0o7BY4r1u
h0TyXmoVFcYznsqfEdtREkqDmxxkfYGTjiIJPyeip9LyUmWLausH7hv5lxu6f0QwtC18CF0Igh3Y
3dbRC6QgtcOHA9tO59luzlsppvz1CRxkywp0VqAVo1H39P1FOOZ11Rh74Q/337H10WjkBbOYzCV5
wVPKSd+/rGE2qRxTMPB33cxKsfeqkLwZNcYx1XDxrxpRU2eTTXwGg7kezHasddusCwe5vAG9TGN1
C2wX3JS0fflVtbOw4zA8qy4sg9TVqjqxj0hjYG2qCn9qQZxw6ZiITjbcOWqyXtaaf33jAH/yJuia
sPi+Bd2p2tYF0h/g5LPdD2jK5fzioQpOhZq6w3Ch6JZE3VcvkA4d1P1JLzAKuStVEWdHQaK+EcAd
mHct36J6TUKeNgZFbkHw+R6xEF29Eq2gBjhN3UNwaINVPgGYQblquPKtV62nS6+eOSZbBigV5cbU
CNHNGsWMsg/fIqacspPuyspbQA+/+tI9akyqLp93Vd3px7YEBg5E16tL8Q56VTCJrFhinBLDIMZZ
Ug/M6Uzhta2GUaduD/JAfpXZc0WSdYNKQfhRc799wNprFH4UbOduvjslCoGcWsmKArg/ISmdKsfx
2hp3/oL+SQjolgwaDHhRyrLw+otCQAUmcbWxsaOJCOoxWPftEJ8DdYq/HhOZ+aqcqi1Mlk2AsIks
0koWpyZD9mBsDWGeEseYveLPGBqAuJ9g15+HnsoD9Uo7UH/k37+hMxx2meoGXxqAEiosgcXXlGH1
DxyA9oXIXRdl+Fnoe+gCAUO3FJUse08mo/w4h80JNfbF6M9+U5v52sHQtoxHkzmospnO2f8pFQ/3
LiOJejqxgq++sn95+zrc83UStBGPyM0Ioi7yyxA0kmLSdKpF5wnQx1qbqDlzyt1ShcFL65mh0927
pc0ATL9K0Xcn0rX8lgge0PZ0Wtwo4InzCrx041ws5f0N6exVq6ptfoVv9ogLnnDl0XcFEq60dYbs
Vzal/ekUGBw9kwFl05e0UbglPw+6kpJV2rjvNXw0yBqyJGGbk2sTVbpYuwlLcGgXvUQpRaxbluMw
0iIFERwrrESqte+PTevwzqnYMI0nAGsK1SY/2vs1x9njjHosOO4Nm/PLhPYVRMumr9SYXP/GF7EL
tIlDHxAS3wb6fj3+urhTNw3BqW/F05iSbb0N3kwUHPKR4A0aON+gpyc6ROJw3RPoas/c4H55U+ga
6Ul6hQf+3CptoLWblxbdX2rztrNYxZS5tlI6MNSKcmiLAPcxOyYyPFbUmheKKV2pKX8G6P8n124R
SJTS7XoYyqXIhdYOEIESYL/PQErFoA1LzsVCE04m+lQionV1lm7sqtlLXOsUTGyCMZZz/543izSE
rega1/o6PBEyF1IE8WFhh+Ysu8fGDO6RpWSJGENor9UUXc5KxqBAK6DJfwM6TJ1/NpMfU11dY4kh
xNbJvw27Z+kumTW3uOh5odHRBu82zOvpOSi18WyB2Ft3Gwa/jMEoRb4gxYi+tueB6Ybo1FploEaA
iEzIXdfA280FAprSRHCzIPHWVUgLz00Vi8uhgKq2Awwr5eRrQFCT//nb7K3UvvJvM2+8yGRS7n7I
+57dgzJCXKg3Qq/LnPzEe8tu8PJpbxjzbx82ya3QKHmhmebUFetLLGJankyQDrWTYBXVv3EGih+v
tXdmYgoRjeHJ+cdQHEFOkqihoLj7C4RoHmZ1D8TRzJdkYfq0844jcm2ZGfZm/yflfU3UqZbtwQZK
zXjlfYAD0ug192vCmaPJmPw9WiBtLT3ZHcPsmXyqQls6ylaaEKhLhixGiyl7JdwlvU2qqT0/BjUg
NH8sgGK+tYGrJcjnOq9emfcrEjDbl21N3SmCKnDKNs3ATyxM/Ni7iH7HbkkEeUMdKOzMCfaxhbZH
cF+GzHD0ZLAR6V32AFxjgSkgb8HwXWBeM7+JHC3Ntm7xiMpd87+ihgePXcV1qFo0wON/N4lmg75M
cd/JNoYzXkQJwMR0/qJI/JkvP03HR1cjOGn1DpVdHig0P4HCSn3+V63clNwx5XoioA/RykE97Vjh
OnsLS2gKP39KptW0ZlQt64WEvnrCtqs1oa1FTEb1RA5me2ICZHqTqfk3QQ2JqYYy9Whe7s9FqB+4
f+7Jujcv18aOGGjFZuPOgsfQ+Y6XOTys8J59emgWHWMtN9EnzleuaAdxmXljlNWVTRh00hZDibPX
QuLSrmgac/VeoSdcfe4C6fZfVoRgB2VpTfz0cvH58CyqmcUBenyOzQWfmZduxcWwOlne9K1sApEg
7eu3VCO2SZwO3cxWs5vXP5wQgnKg0PiXB0bVk8eJjR7ZpU9rqRZlglvGjgNvyau0motudjFhX0/H
UYyfGoTV4zkgk44PbF0BhXJ5XrrBnD3hmPkvkkVaLa2Psi97QzLnI+TVJV3i1dx6PzNZiNa4x8wg
rTqJPtNtoeZ/tDtdgHXpPhsKEeAlJhk55QUo2WX9OBHSFoVf+vWDj9AcyfXsn0AKMxb0eMGnxEbB
j14MBj0hTdbRCIRn4b/+CMz5CtkN7AE/XhJQtVcV7C5u4KrmZyaXbpdVj7zn3h+lT2ms4ErfhMnR
J76cJgatfUES5LMqwyIcaVowoCkHawrkIvDqH3Znn66QBg+0oqnNBKerUaG8sqVvReN5Im+Uo/3L
+UAFRTj225v4xGBIpiZzLyUhEhvxeehlKrrIIFPp2nU9k7PfwHtypRXMwWhaBSqBC+x+VhJ1U5Hm
ggw3U1HlKkcR5CTz9dEEjPJWfX7OVB58YHIwEWkJKchYCw+sVJiQb2kSUOMOCw0Wb92mbMELICGb
B2VmrdXvWjP/B0Uv1SbDPsJIVNoQkzrSJeQ/ct/NS45JJXyVocU2Bw7RU+gPWxnfZws7xE7+pueb
YkQ1yRVFQxPy4L+Inee5EDCxT3lozFFLM8JB1hqYcMfBxqZg4e90DhmvIbo+FjKyJH4+B3wCIt7K
X6oLilP54gRS6Tu+GFb6kNhFkDYXGU+lWLV1d15nweywBcp2Eg6fF8odopU4D14pV1CSF2Ujbr4H
9F+eg8b+ZpkwvuULhOFoEl2hsGoyN01PEOg0JS7QJMD3EvXd7SfMUVYUqX0tl4pd8oiwSTcoIbqs
FY0ENNTBdeWfqR6uyMRbqzKMhIGAfW6Q+itPGXoxaA2MaSWYSSr372C3Erp7CLYf9H6o6F8Wba+u
a0lOdzWcqHv4h4FkRt1vEVKt56fSnDGQVJi+e8dY1mC8im8yGN+iLsKoU1bDGE2jzjci+DWFVdjq
LKLEy6L8bpBS7UvwSfyPjQvNnc5sivR2AS8axeeo/yi5tstlcVG1bi3dvfsS5EHycnBV6M4xrzD8
idGF5uJTkG8jFRojha/BMXXvq666n44kNAJEDgfD3b1HW+tjWnpWQakxTc9JViHg0AV4b/xx6HcP
Jp6Wf/GKGWGm7cj4Jw2Oe8BAXhnwQpArqLcMp5rMFudDEe+pPqiTWeo3MyGQ9G2/DrGAjjZMEMn3
vOnqn3edTt6bA58WiyFUcxB82dG9T83JMt9Au4Qz+WKPD++nzn0hWgXIzuku9dCK7IVig2uvP95q
JqINxgKxJbM0nCOL70rVbNZH5mPUEXGhWJfv4dRETw/U4mlHzYb13d6bk5F68Q6Y1VwlPwDaU2aH
GLOgov79HXB/GJH8Q/9U8F+mZmCcKCdgGIv9XqFLjG3cRqU9MH19lK0zCjTL/lejBPYBtXtMKBQV
pLLKnbqRcnEq3z2R2WN1Ny+8QbWxLc73BKpdWrSpp6N7HVPLb6woVo+RoaX+S5QogarOVxw+wi49
za63b2VlVIvuhPL9IZV1DxCdKwBfhi1iUpdaIFFaGTNyZfANIzo4tVgDGRGaAmwkiCin2EH9SgtP
rOe1zdUPzlmrnime5yplvzP69FQ0mrQ4nC8mAbEUlMyAUan1A/YvFB/7DjphFcHqC1LBjS7x0QIf
VkryRgCqJC7I6N10U18RO/B72tYNI6eejdicz4jmjZGS5upJ9/I46A6ANHM3M6sDrXJe0cQimzm1
0EumKS7Cv9RZvXFY6Jl6+uozw0RnqbSnv4y9HS4GQqGMtrV83N16+pSpZiYw4RHE+QthurMMFZXX
GCIBuKY4nztg9PfK5rsgok90XzgNZOBr+97QPpucoW4bcS6fnOhB7dH+h9RuNpV7TkyqeOSYXY9p
Ce+0Eaw0W+A8AN0P0vVrDbulbn77Npc78WVk7GOanBIbM/o4CJiOdQFducGlih9NaTDycWyauFq2
C+UKDL7aR6IYWFSWeNFeb2VFI/wp9khYjZLG7Ck/mA2hSlkYh/VbaHCT5Mz8+1oEm3StVsCAhBHr
QQ8vm3zCjsFpQYy9/VWbvX39ct6nGHJ5nGXrfPm4760cmYsUH9LisFmrnwzofOuPMRi2eAlq5lBk
6vU57mQMzTqixiDgR5/vno9v+Q6/q7QZ913rQPUl/PuMupGMey6XwhL8VOcXCjWTz7B4k6E9Z4bx
e8LH1YZc5elhPmozjpUoxVWUE5FsUw8qjzGudhLTKVWYoVuWmWJj5RpBHDJN4QHoVUwwhCvpa03P
PR1x2Ya94ANCr1/1fPWt1FP1mkUuQcnXv0OoG4LxMFgZ+NvluyvarsZide3SfixpW35nxaKvU4RB
qGxyFaLMm10v4jb/gcpgPHEu9IYYTkumGWX2XfpkkDv3sIBrBN7dNiklTeXeILaBmYF4bamnY26u
GZfmsL8zyLl1AtKqtT7HZMDCKxfPrhJFdPevt7tnK3mZAe9C12a4m5MXMM/HM/yg7eIJ1BFITYIA
oNTVDKJy/z2V2brOjxjqtkeCvVdxW1ISwmh6ZyW2vAlVEPTIOwsHtfr1/Xzm7DQrFfO0q3ymcwgW
yI6k73/GiXzFoCAqvaSUia67+0elI46hQ+yiCOrEnv3ql0ioAwfkm51EsNiJHYID4gu5M1Dne3yr
e1jsQ4ec9cQpIfKAXeSAQfnyEeX9bryfrZWa2fVROsV/PviUPJotDWExu5FP0pOPgRl90q1DlMtJ
nxOvsUmym+ybblAUamsZ/oQJEP7PT75ZEA1ztmepE4YVSsm7f6DyzczM34qG7/Keb5NYhD42+jLd
AsACh1I4mkNiI3S+fmm1SA6zJC9nJUB5PW6X5usNUSQRn5IHgu/VWCUXr9TqDren2K9I3RHDO4Zx
vjAj61sJpNSrRe3OpmOPBryeeBlPlqvKcB3zKI0zlEltvSisAVhNmxm4me+ZAp9DxgMZildHp013
Z/5wwfI2xyMq7QFnimdQ6iCiw+uwmCI5zpFswPJRIrLseosFViy+6573l+WnjS9/MW6VbdxpI4JW
2UaM8db6L44IYqcuYGafXtAQL7JvT5ryIgAAPy3wjUQOcUMKXJXkb3ErG0oclQp9yIASEQmOsZDl
DrJ1j8tkA4JAfSGKbAxjBNSBTNDWZJm88JROYPZ9/caqmcRjJqId2BKXn8oxRQirCt9a7jZ05pve
WO6R1JPSyJWJZcNqYnCP0GsiFKqppGtdeeVnL3AzcMhyh05Y0I/U0cPcoRN9ygJpCyUysn6yhXse
HLrNKFbqFtT+q5cLpgcL0eDBIOc2gpUAznPGaeRsbLNlhWu75XS45dqqOaHV9LyoInC/omEPbziv
sYrZ47vRqWK0BWP+zQ+cqO1VHtEu+FA1Ez6jS93LcrY0fnzCxwZCwpDSQrfpzuHeuNUOvauEtHLs
pH5mECLbxk1vxZfJlMPcN7u76QjbQRy3bea+Rw3PtxpZZAFOZXI4rtFJ6OpC454QJo7YLD8SrttZ
TYvgRvGO6mhZDFpkaG4BvhvVC8MoIBY9Xs2a9MlEm/5QJF1erGSI+dPuplz9x95O2Zu2iXxp9LBZ
w4QnCDf1CrPd+ggR9vHHm4eMv7rL+CV/ZCxm22eiDEjNSwYxPBzbcTMmxURezjd1C6pah8DOIG4K
GBKVPmuqqlvaoGb1TQgfcGy8LWfICi6SDx0G+xUp+3t0WxCvXix99o7C6DwI4gLt2tzNJ1zgLkJB
Y5t5vnVZsmSqicXGi02lmbWwBouss8rPQ44vSAL4ItvJsjBpapa7CuCipCBSs+HGOVwyREarUNQY
kHjmN/X98ONWJq7aGZiZbblLuF5VLY/SMOdfu7hBMg6VD6tfEwBnWeJzl6XIqufRxegGjwyoAIWh
kNcYtd5nWj9jTY3Mooh9l4JNTWwZ8beSyvsinPgM/hM58/peDAuRJRJh3IRoKaPHJm9YO62SN/cx
U8wMY7ZtCQmqvAZDE+8M7OoucIY5XlNKlyYnFyU/aspAb+uVXadUzbhD6h16FwpMpe23cdDhZBWK
5rAytkh3s+BiL3agVxAHroq2FJBsWH1Svd4OWHnCLmKidJxTPTIwLNXe5ndWQRV/O8S2pbvvwshC
L4Vhe9RuzoWuL1i85rvXTSEc8ftkw2rT6n7eWO26lou/b/9vafBv7+amW+4eHajYyXVXQsKhgGBv
umq8w5BfnsGImlwFXuu9u3D2nS+daTSuTOJUfmBXC8XL0c+oPCt9pWNyNnr27H3CiT+DKHvZLECG
hZSGaW4HPgZH/69L9MxIm3WZx4p3WLLLDNUMGO0F8Qh8qNKM3Nax1VeoNu0uo4vE7ifRvQsvbZsJ
EF2A9Vg+IA3O4MfnQG8x6WESwaUA9YUwYR+HXHVMUF2BSjol59tUE6PjI5/sdXI7fCEV6E7x+iEf
zEs5i57AkS1bK5MGzeAFywjmJ3RKA6h38lZOf1F9Ort3izvQ0M7/tnDjhl1NI5ezjEDikWHnN1wv
eTuAxYKmtQRiilsmiqEJ6NCs822MnQlpP8EsW+gehp8uXA1HcKHy5Hj0osjfyqd8PeZ+DzM57NSB
7poD6r2sUd1yzaZgCULGEfomi+e4WKn5FsZOJkhn0+1d7nESNPsdYcyNf32gR1bCfoTMshvoJ2wg
IFWe278YH8stwW3a3BAcgn3HD4DottPrg1YmJT5APjyy4A5W/Ru3zbSlO/rIjFppsOM9bc3Pucn3
+UT8gu5n3c6aH83pORna0IveF6BCnErRD8+8B2Yok1SeElTOI49lZ/81zN/Xq2OFef68YEhnAyw1
7i20WahP01sIA6QGZSWK4NI2ugDlutK7GgaJ2SRaM+mG+aVUjHBvpjVP6wB+0DiCQewOw33VVYc7
V9adT5x6yf7B1as6adtOK34H7E1ka6sdlSDsg2rR1OZWSwEENRm0+N2OUIwSZ6tFDj+fAQkYHaia
pTbJy7ygRirtwoZMaYUJTuX/qwuoFzW/50k/TyP0qjiRGYUrK53tIyV5bPiKMvpZWbMStWBYUim5
Bex2bBPj4pcXnA9IPHxKthX0VcTm3QPcjFomJgJ9zpsQmizz/wvJnSUef/eNA6J8vLUxf4G2bgC3
ipDG/+pOTsUeiaonqcr3q8MJYaA+YuyuhF28VxZBntjrrsY0eEuHJBP3VhKzen9+E33e3k0j+ZPi
aZDvCM4fvHQXPnPW1RFIcyK2VweyTcD3S/G+2wnIjUfDNH2X9RNDI0HaLUM/QMg3SkPGocxZ9vht
Oto3k+IlNKPBwErZKVwJ1tIMvnzcWmxlEJecMTM2oFhsXhrQIuGaQRzrluzm1x0gLlWtygDDIj1F
vUyXoYdAg4+rjEbpMNqsuLhU0Wftbyz7UVv8TXj6fe3GU0xjR3hPgZfp/Ka6kAgK1NvWNGuhR9/e
lJn+VI3psrAiXn5zjGGsDptmJHChwjK9kvuRHEWHWEhTgbzMzR9fMEuXO0UDr36n7vAjWsDMS22A
0xlGdPt3qvP7RjklWV+W0S86syNTdydG27GwDG/UyD9VUPtMpzEAZH/5VCyWKWhn9N3MKHrdkei5
fv1WlBHHlfowrQ7RBsedp8deC4vs7f5GdylMlLRlM734o6ageKmz8vH9btt/0twNuNggXi2DEQ3Z
VPQYexD/5junuZ4uxpZPw6akt+VdBJBAXB0SlrLECpCHvFmJgh2eD/gqUqndVO/JmvFgG9Uh0kdV
kiCzj1FC4d4Fq7Hw91lS+7Cx56Cna35Ksd5mKL0IoM0wlZoxjbI2uwTzlLKtSgkcRwrZk0T+zSiW
0iEcxmNQeXJQlIcPjmj4QEOANqKkFDwdJfUnVRDs2rjnaOg0CRyhRlpqnZNgbXyU44WHQEHgzJ2w
yyndPkhCnU45yuIwaIo3PC85GbTieTUKZM6HSInFKwvGJS+CvrDJxJzmeRb7+EyeZEDVsqlbfoRz
vEh7EcHCv3ykf7BUIfCUhDmL6kbfdJXphDz8PdoPNNbqODeZzMGwmF7pFWq/LZ1RQf1hkVNhww9f
vQEbS7gG47qtS3KRahf/QteYA179RS3rDDJ4iwTVYKLvCY1aSYI9YY29xaHo+pSdnnW3eEVirXTe
KTIxQff3apUn7H6Xghip3oXRWKD4rr8xeFmxPiBPwOlxIEbA5M6AxgyvXY9L5eK5C74Gpx+80fLl
5meHqH+m7rk+zhnrb+2elrMmyM8+4qhnfuyEPiFpndYKTDBQGONGim3tdiweUxv/yzlvDq2JOQ0P
G2INrIv+ftkyx8ZRqybfgefR7W5v2WuyMwlhyYrji/XS6fnBteAUqQg4k4UtK1Mc4BcJAhGuWJIn
38DmqD06PHIz5zrAW7PeO7ABUXXVEhkrLt7dR42lDoBzBkuAq864TvP9sVKBqCJl/uDfLVJwV2RG
bO110f5krOwNhtx+Zye8Nm47JV1Ms6q46n40sFOZeQLxET2w1jvr9/7BuOjaaGNmQVHbebJ5Ufen
sHvtW1/d1K8G1RLrDmu7hEO4hpLgE7gAEcORGTWSTJiUMF6kOyGQjroCgAaPz6jb+GDTc7Nh0Owg
wJLMwlQhEN+qQszfTIMcTA3H7nxIOizPvjwSmH5PJ2Fy5NzbTmHSlT7rntB1C6dOvaQe43wnn5tX
DMBmvQBpaD36nfMABmT72T5MamUQaQOI0LLk8nW7gNE+AvrTgrhL+eCrDTrkIvZoTPVhPdqamagr
GZdxHrvPK0yiSCj1paGzTOJIDNjEPJCwDVOwpPjfN1mUp/6s2shWumcXPDHP5sNuAIFb6MSRMEAG
QJLAhSRABG5xKqB1YcJ6pUcT/LAibLx/U59ERdLavym8zVjbah6YqGqpoZSNyVFcPF6u34Q8uLpw
BohV2P5yOWqmhg7QqNO5jQMcy4JFyUS1YrQdp5xntveK3gH2grfv3fp8/EXg4YHtfWGJ7D+jRFPR
7Hu6CqcPHDjPWRUWbXN8O8RGldsm3WsazpZ7vn6QmNa8tDNm1SemAUklQUacf4cUwMzA8lSR0xBe
sa5WGpjgwnFxS51Dlwf6w98wlS8O1bwV6L6r+O3L/PQBHZm/SELiVfg4soPDyN9LTGInWnE02IG0
zawN8ReM1rjklIyOUnLxIE5o0IO+vvDiSu5Ppmbw8h0em69im8tlsBRvLkwiWWKU35dZLszHSH7r
2Fp8lmRwf2ldwFxludMsMbCYD0Z0BrTceivLyc3wKvc1ktCcjIAmXErpL9b6Zu2v5u2zn6AqskiQ
JHomcR7syay7xys78ez/pi7YpVlFrG3UqxIjz6heCVEZ1Ouk/zGLSZMkLS70AFZKy3UMa0JduZMY
SFEpX+OkZPXbfLU6/SISnZPcQTpNsxEnL+hDGmwK8tnJ/PUdPM22qtJFrsmLq6dzIvozfCNX4faM
3XwVy3zNkmxc42190wMvAmpWS4HWwRzlcM5MtTFInuniNrIW4IANjwWoyObsYLa7LwZvyM3kEisb
FK6Sh/KZi/SGaklH8Y9TQwp69FMK/9nGicjBQrd1x4b1W5L/qf+wd5kC2Ghg3mSoFFtRiFRzMWUo
0Vm2vdKcdazWsm1imFOfTVQNyx70jLRGsvHUDb0ZwcXKDENqeqKQJpd7ZyrIZou8+pZOlgIIyUHu
oc0VicGOCX2IEpbhn/k1kpAq4mhcvnA9EDGY0WmJviMlD/GCSVm3C9PAfQDlNXMbD5mzRixuKm4N
gBF/wjeawRtn4Oo9QIGvymCwZQ5+YpvSge/8QQBLHEUyl67B1GnNI3ilsGe0EW68AshW12nAh50V
0LOOdZzR2UsFdfvNoJhB/3xzSFJD6uhjs+9+psJ8UmzmP/HPoFWPpwVlQAYf5RcawHB46KZ24Es/
todVoFmEg9qA3VYkSpTkvYRDiAxulaxgnLOwYUpGJsepW8tLPx3jK9hDgn4xfl2klC0NKy1UOvAO
BbQrvhaw/rBYmhJFY/aRz8sp6jyrL9DRZ518h/CTkZt7FtTIqWPk6wTkcTIm+MTgMw/UksYa/B5U
0pvVk2kb+vSzcpXIB4m4PteQ5RcLVVhSRKP7tDl70KYSagiUpi1z+hs1qkvaTgFSkNI3qih/hR56
Kw/Et/q6QKJ6NX/DHx86KRRjBMdfFaqyJ/vxs5Qi0MQX//Jfo/dLuomiPPkKqjV7vHSjVFs6CHQe
i36AAUTRmK/0kOePXh9lpMP+Js5PFFgWqjrVlEhoknK1hgvLYY7SkR9Zk7keEaQlScn0P6k89SRY
UuQG/sbFaflHrMLLHrLNjPwr4aqQ2rgNigFkybfuBPTfaK/Pq4FFiHeawgNG3sQQyQcVa+Iorc4K
v3VgA6xWbH/fQrxGfGTwf3DFPSa8POW6iHdTxwDfQdUmj1uGhiC25hrxvdTZ0GF2eIzip8BPPK5D
6ga9lTEF3qzNJg9xh8OmtMLA5FP16CQvrqMkxq/V3vSbQA1XGq2z2NJbGbNEFQItcK9u1LhyKE8e
4/KpzrleJxRI6aiRFG+J6dDobjCu/rWbOoO+O1p19vfPU4bHitjuMhATeIlFcK4OZ+aQUdgo21+q
ZEDTvaMPXKNTCptOzfs06+VO/CfZZfaMAnjpp9hxWhcuth1sSJSMlBjqJrOQ73eQ0s64bxSTaK8V
dLOMRZ9K3ICxEeapkeIxpH1E3jvts5IpIGeuUW5rZePzjZrfAf6oL3eqCxLBTSqeVo3WJ3/1ZugT
VpJfZwsKpU6N8asdJRCnJWLHWk/BEH7If67uY5Nm/QTjnaioklwUYNR8eGZw6qNJ2VZXOvL8eqpu
KjHO6IThrMrIDmRjNoN1d99SapJsV90rZeK9lG0upKx0OAWB6Fiwjkzj3nem6AHovaMAaVoOkkP+
oWizrHH6cTTQqEt9M4uDk5IpuC3+/P49tRS4gjkmC8yP5NnejHm2pPOW2kSBCgrb12TbuahsENVU
8P+WuvLwHpZXnTXg6ndtcnC4ccy/32GMDHcKJ2FeSYF45hE79my2FpVbODP+sVvj2M2OiAo9S/Rb
VO02VwAAMBv7P+jtMOwOrsL+Y12yVTUd7YoQOq9SRkpnn9eofwijOOEldmMLon+Qq+KWwGEwEmgo
b6g0366iNxAvaqjznHNNO2Rbe3lEIERVC2xxyZqEATgKYJavxNZ1l61NatVbq0mtv8nFJC6QXBdt
BqARa35uOw7RDeLFyzZ2EyzJf9joeRKnWRNfF8SoSxs28ch59UlT+iPrkG7dt45EUzlK2ct+84ks
Xjr7rir/HcX0CXOrF157JRVNtQAgrHFxd0xngZtnP53RbZiY7dFtc8+PXIu7qMAKEWDjmPFf0M+O
komFepeX57bZ6XYFZi+H1prM/Oa/hgfn+sXxUbz+2OMULOosulVV2n4g5UzUkZosycl55R0bmLJL
Pz2wjzdrSLu6vTiD9AMR6ZFTvAKI0NuDEuGxIQMw6y15VgTie99UBhXxs9l10iJ+ao5IgzDx8K46
L46SRdjA0LKvMiF4Q8WY6rY4wWkRc0t8CQq+2sWju0OGr9N6wi0MRL+WFIqFJtUBJQZF9bJJV0dl
u3ZGirNCwI4TeVudUhdfRCtskPAWS39kR4NOMt93MyxV/gdX+CwxRmm7OairbKa363prDL3vmZpV
nJDaNqJFF/tx37szKPV+asHdYbfZ0lSjlcUegaHW590I8QwdKRxnAo9iT+uNWdxhXdK7sCVl0Pyl
i88EePPCbbHg6a8DuIBiNmGS8aAo0CYCzSokY4SdCfK2Jxfp1b+7ueaqKEYG8h04uRLN17MHwWDf
KZukEsnK3nMI28B0YrLMUgqSb/4vtB5O7ZcXYnHwQu2IXoyku0IoJ+vHTCn2oxH9pfjokd9Mj4tB
zRirCfx+EzzAGmcu0aHVR51MPfncm0PlecK0NXSJCXjTQWy2vSv2wdWgIdDE5hU2g93k4YeIvENM
t5O0+LgriUXnvA5AHdgcg9O7Bj3e6mLUXrM7olskmSAZydaPtyC+y6a80yNmh3zAzirMXY2yU/Sn
nBgsTPcvk2xJcZudlHBmRkZrSGE44cI996onSCMUqCJTOrJDd1t2o+Lke/etAbuRD/2hWz59ntOy
raw9CMojjGoS0INWcHb8tKoNvVX8al+y/ytrlk2M2hXnGoC7z7lS4ymmVdxzIbAS78mAlU9N+Fzq
zKX8QV1RkFqw8yMmdoH5JhlSWmuBeG7DwWG++byBorc+mduu0VQWg01dgtGKXRUXHhZ7VXE0SozY
Q3l/uBz9k/tBTs5tkMsv0HOxZLZ5RjAq7+PM/88HF4/hlaJhnImykbwbQCfZU8C1PFLExIimnTHZ
1zskez9S1qoPIhI+TV5jnz2AFVGhCQRR1QixbFOfbV7mA45tzGhumSveVAbHq+FA+xH0tiEj7t1B
jARBrSeW7BBEn80V4LlEQgEsmyTWW+/Fg+nxxERh+IzrxWzRTIfcs0fL85VEQTgLASIl7q3ljGLP
oR+XJkeaXN+bJESZNOjfVCK1mzXr7TN+IMFUoJaMMOjii0tj8E/uF4Jf8RhjwphaF/iXHeyf4ouF
ucZjdli6elShCaUsemqXPn1UOz/Z2E8mE9b1BH1vRco6YeJFaIn+upoU3PPF1k0N7KKnECGrxnWX
5e/i5985WRtpmJpo9uQAHgn+Xq/zkdeX4UDZJlwklzy/7tUdTaFHfZgy+9MJEzaMGPh7STGk9cYU
kMqRjoRYvsO6wS8AAZVYV/LfDgxA4lWdzXbMUytchsiO7KWF1Gg4BxGH6s3Vb0I1lxjKjq5F4Ph3
ROVFpV9WNy4gYZDOln7w0BcW7wi8iQHIVrPGX9/g73tnh4xtxmkwSUBmk4WD3DrHKFHPONEIBuFd
S9j4fCNqplDAhBPwv/jauaCsfyU/aqZ8udEIqJRC8FUOgyJXHWqxZ4WM/vwCzYnGHTIMMu0A6qOl
LrKZ2u1A6mR584prGTV4oqO685iIzgQwZRpptoDSVMLqvfZA5ajDX2/2x6Ap8OVeOWeFfjsi2/xE
uI8illRWcOrAnInXgxQqWQzi30Wvu2JqRF01Igks/pWT7OY0V9w4oYcbenJtSyJSjvPjuk86azpr
1dg0c249gtU+ZRMc8Pfc6IgtwaWb1n2qLzDk9vbYFztJEx2lNjtfoncItL+oFcukn21Sg4DMLW4w
6xv9RUTkYdrpXm0xaoIBcXflXIeX3RimrxL//Ts0AtwMKv8dzvFqaQW+CcrtREqb/vZC2ssqY/N5
bfa6UvUywKt5K5pvx71krQyFRVpKn5x119NW0q9yGgQiznK0L5mCUR8qSaUeuFsH63mZTe3Ztmx7
abv5o1zfszlO1lm0kWcjbxoykXe4RH6tClNSOm83BLrQSIea+HP/CogrEQBTK3sChViNV7SsvjWC
Hu07zGke/g/WPCNAtvOWihRgjfpgzrFJ/LaBEszVPWZOaUvJFKCf3w78rTv4G7geuG9tuQ1YlcfA
2CLLhjTtL+V/IkLHKdn3QS0Ktbwqh94DHPNlBHNV92VGn9qam04Z8tqIUuyOUHGpzpl60DmvZEYo
aBMbF53m5LTVWjBykQy+6+6UFsHAiCvDmlu8KSWyy16UMG1uWn2LRCN1HGH6Z+9DUX515B8x+389
0Bj1xJXJPY3/mCw5WufIC412wDb7XCruVkZmzq16jznoJmeSEMaxUurU40pUhZ1w/lUzdAOH2R/M
QYAZJvODrgX4doIAy8aBIU+Sj2CJdsLK15sfBvk7voyckOb2Ht2uYiy7cQqeJaeEsQt/YBMtTeb+
akp0mpVmKpxIu3WbiPLr25vcTQcqkufXgzzFyZdoKR0TyiW+v7GHGGJ2feyVeZQZk8AZdvx58KFy
b0RxBbavGsCpTqHtCLtFRygyJgGERYUiCmd5Ls7Ta8DA7QeN3CY8ihqOArmX7Lt6X6qTt++mvI/X
N6gyJmjUlDrcxKl7IiG9oT7kKrxTquerPJ5XYdi4is4dibPSSW3UbOz9fuATd+OK7R1/wBKxn5rI
Dithegpm2fc3I3dRuzRvanrvQk02YQXydF+wDW/CQiFX7RVugMIJnq34aUj2tYkFV10m8kOkYuuR
COdE3Lzp+XppWjfjLYbf263EO4N5VaWHz04+UJ32WomjleHAfCqK44H+0Sz+g8UJ8aXA3G74PvxA
GjsspvQA8G3h7jDe4+h0+9g+vUQh6bCogXG4Hbzyv8E+55A11i/M74H9n84dF30Axut03vuVnvJ5
PpMie1ZXLUUtEYCroiqfmEe2m8VYa2kXYPVsYJbVf4yczGJBEZSqOK5IjRqKl6pH+wd2xjRK0LVy
/1jfCpVN+Vpgi+7jRt96j/LD7PVQZRIDdVGwra/Y0tkAmAstAwDIgPX1CWzsBiHZ1osIHYV9nsLN
1EQZrQS7p5NYSqInJAKEIC48z+oxIfhpEQp4gZT11kqt7gVIddiOlsVitNTko/1uzWY0DeNJmXOM
+O8hgVyIkt9kSm26AGCfMOYbsQHVDjdURdJaeZDJOGw/nv9BdXCdWKneB34O3YmoMnKM3NToCudm
b5uX2rat2GtPfV7M3X4LwdGvb1uachD8i1eT0gP0F6zn5BcfQ9taVYn4sRsYAmQyK6UOvsWXcqIR
bAB4YeYF1xlQ0yQXUoii3COUjsYDvyXWi+xBnN2MSf1EWYTHq34tfHnI6SdRrRqoNpKqEhooZOmI
boOiuXFpb3rzPyMGPxjUpZf4weuvvLOCoFtzTFEiKKYoTkm888BI3PeyeT+JFM42Kf640i09PruM
+PislO02mQXOdNAXKgHmMz464YvR+uvPPCfr4mwgIg4mRdn7soS7aHmlme7kHe8DSzCUeKV+xhRf
pgxeuEMXhOApu7iMnZkO64nnfIJARYnimR0bUPyg02UPxznEPX9iPwkqaw2/af/OP4M3V2W7oXON
weF9Zv+KuVQzVxZyruIFmE/Q5G/DpVOLp+7XnSnrB8BmjHrW0+aiGYLVGMkG7MAPNBix6TKwTP0M
NBkiGKcF0XUqynkLTbDzGk2xnom3FQUnlCbT2eUXvkY6qnf0HYUC8DhOCuJFjkXM2UZG2v0b/RXc
Aay8RbzJ6LQqVbYOo6NPKbj7WBbrOTyfBFUcEICgyTEj094/BPKVEWEcaISHGl9StWW0l4A0SsXC
XNISqnjWZtw7d2rWdTOyP9L5ix6AcZ0VaOj7++cmi7xApkaD7HQ/u+SOQqGEAzPiSuvu1wCLoQPC
TE3gUVaKwyiq5dqWVpal35kun+YIaLUb3xoilo2B7pMP828XgM+EEp6M0qZSHMQCSTFLnU6qTlJC
62d9sm5yDVZsYEyoZjgFpWLMpoaimQlD8gKfhsHonqPQMelAhiRYrhwe+W2wvNQ80lkAsJ7zAwQ7
mjSNzqlo8+cWGvp6iwfelNnN0LNizwWplfJPkj9mta5DdwtOF6/8/k1+ce7pYvnXErKUvzusbChb
MQtDLNDMQ0vCcy9p83IHmWVzm8IIrVR8t3KSNEZvJt8HtafZ8U1x4950lJwmpmguq5pW9qqeM1ry
bPSTMw91nc4zZTDVym+qvKaUET1dggk6t3r/A/XGur3+j3et4nOOfm5y3jjaEubTkT5jQxpGXXRd
SxPNcxcUR4K/iktHA4v0d5GSWOSrtKNzpAknQWzVtPsNYJ/pQMELwS3gEgESoLRV2EeFvk92Z/F4
fPr6pYwaiEDMenol2aHc6/NyK0s9Phb5GoB/m7UVaNPE5Q9drQkFOlP30n7sj9n4wzcB0KwE/2YR
Vj2OynCpZkidV9WJHU+L0IhOPLl+X+wdeuAIzIMkJ9Io/giP30bWaeaMGt8IPQzjnhCtSjHmZQ4w
6kMye+RkrdJkLFFiT2r0K5PQtGiFp2P2/0g7ZLpNftUiUqaL3m6juWMXt6HvAlD8v7l1wzK5/tcZ
8OwCLfXpWXtTviGzyzTpjKwJgecA0n8rIfjiCoRrt0Rb8fMOoGcl8C0XtNNA1T9hgC4f0odlpbYF
ARExmKM11MCf2Vonmu2SEqU9roiTb+bWR3vDDCFmIcQiswOL8HXvcEIn38JHv58aqpl0Mqq09njO
6Z7TnOd3g7Y0fmVrQqhZo2vKqcRfanCrjakR38hVJCXv9v60nzydrcRCXd7dey8iYMqGtEG2nig/
PIOuKj6meSFEHDitDWadIpYkcHI0C49Vu2h+y1Ue5q4gK7z2UJJ6QctEaghe35/GOL9EZBAbHi2u
l75Dp/8/n5p4fJCMMIHgF2O0TjTdFM0XOinqoL6FoT1vJxs7JR/gKON4OrJQiFb1O+6qN4MmRUMS
Q98+ous5Cp18gO9HA1l9vr1KAVW5MQemUAcro7AJZLCwE0BhE833SwISwMWZCGOqL77d97tt4zk8
rJDpFUd8lKRcadmyxuW2oJ0Db6akKROFEjBoA09lznbC7qAZ22vJhd6xzh+9lndN7DqfKzOnzBfn
OKFxBfZ4qDhz9jb6vDozoaNGdyPKLpS57To/FiyPxOmrXCH0eRPZvXWI4gtl6bCKw7cSSnWpqccd
8YSnR7VdALiAf+unKs6JXPJMCXg89SMaFkBPwwil1rPMJOmrzMj7igwVyOBs/PHafSw61fXWa3sT
4uvB2/ULa8hw+Jkz5GFbu7uZhqUeMKlspMnd7/eemciJRRGYlHsCnRf7ApsHslsK4rcaxgxXFGeJ
6g51Qc1/OxcVGVXBOdvf4Is98N1I+6QAIQLcKEzlIdE2i2HJlq8NpmxMh4L20TSKnP2Iqb1V6SE7
64SCuFML4vCeuMdr7KKah76c87plBOHKYnu/RTKOv38r/IFg4Y8/FVFLyq4V5IdjNza/dpujtApb
yAO5btgvSYrvZ2z6cj7UGxdekzX5/UQYgze4M7mNYtsPyJ9UX0skzk14ZMyLLNNI/JVqYxhmDBRb
/MQJ/yVHNr0rQjv36/T+0rROrnblpKvMaEdwbocp2TczCJg+9JXU3ceyC9gqCQ0z6fMSE2jjY4dZ
vawmIbYFt7HWleDJodR+5iqTgKhZb+zffB5y3CPZ1xGupeo6++O1McPHSaWducwOCIj+5gak176P
aaE+OnmbevigCQYLgCkebCumjx1n793cYBn9IXU021uPb65tlfS/681WRft2OBRE35UVioFadubU
9+HLQoMmZlNb+/+/fbqIuB/EBlNqv2jUWCK5s1DrahP4Jgq8bQ5hqZeJOKTkYXZHwtwxivplST13
kwnuV+BvXjbDERFajXup2zZ1/n9K1633Qxi16kSLM2XJ6TZH+QlHlA8dQHFkY/D2gre1LU1KPcGW
zxK+0TCRk6NtVDn1xdzPSvhUrvl0+nY4vkPTAINMhHksF028IyhQ+AWRh9Gg6sYBci/O2ajkEQax
EDxu32Vr9QzbdFsaRUN+W0eBNcl5jfDxs5HNEAjFTCHEH+ClBnlmW9M0oeAOtcFgdbVfbiy7UiPk
qkcMyZ/rzIrOnqZ9ulGQPNL84JYWp8mitEqRT/fbhAkYK5acpszC7xEITyhbBYxf/TDPEY8MJIxc
8Jur+vMmhT50DygCecq4EfItqPyBVFoLvWOhzOko1ojtRyrEl3tTpQnqDSO8TNsm4yHcvGl3IftG
61AxaUXBlO1QyK4I/OO5lunp1/2kC9M9Ykm8On+bpEPgQH7oY9JBGFljih4J0uJgQt84k5Hv07Mb
IsTmVxktwO61hYadIBoz0UyNfGn412qevgqiedevPVhVcJwWgRvblqH9Zb/rYCEqvwKtmQon4AMy
NESsgAmV5O/rLZt6cWFHa/kWUyDqMbKSvzAp5+STQ5YdEfYflhNq2Kuj67v2v8C5nBX4eko2z5+f
rXF4096IshF0lM9Di/C2nstcrM0B1ScquJNJv4/1SRjKEFra3VmsKW9LrCNioHHcRGVtaYQ5ZMWb
2jzt+jOaoXFOq3xV5mcA3Q+vioZgtEkwuf9LsgwmO9Nn/AANIPKqKv+D/DIVZyECrhgg6eO0Om+u
rhF8o+G0sKfHBj6S7d2BLqZermqTJ16yCc/ktbbUYVNgVtVqOYvMhOFTNSgamq40FDaHlp44mPhx
U28o2TsHlu4vKJTZSp8UHh3K6G9h4lBNE3vlTM17oURN1NAlZzy1sJT1OzXdEAl6bHnpx1I6dNR4
dB3vrUdJDcq4H2NlyBrr+22gq3aTU6MI7JJHc+mqO+0nQ7DEtBbZbuSzn+I9c9YoWtFJqSMjBGK+
JXRxp8/H+JV0i7s8QYY6wLLthaQbS4fFApUf+b+uSOcZ559gmTv5RmDkVRWKnagqmf28VPRr3/r1
2jZaOF6BsW5NjfuElJKv+jkpoR1NHgWN0qFEzgPqpC6x2918xDQiUQxsZXBfkGHHP8gmbHWocZS1
0YlLjUr8FonzkBE+xVfocH+U9ys4m9n9jXT7HcxLKUk+ZfmehAFXTLSL4cXbj0KveaWxIJyTqrha
o572QDW1dDzYuIbqb3AG0RqD2Kuv3x73PBlrf8UDZSrJMIoDWWyoWK23cGIFV1t9jpO5i92j1wgn
oU+ZVOnAr2tPPuuUwXOASSL3OCTmCC3RowMvspYzIIUpntkDp3+QYtoSB6g5HfgAlUjG7Z9/Naq4
3notEizqwdIv6xnGo6FsxBzMZpx5JsX7kthGU3DYfN70VCG+HhsT7SWQH99Swa+vo+x8hc0ju5oV
K7pYQ8nWJ4mlhDkfDWgpP0O59rwU6ekso04PxFYylqeYzNJCCbuT2nDsmHWlCpjYieXL3HMVisoo
2yPU0VOsQYfEELUu4ZmPf/IMy9ZIOdkQOTyBHNhPIxFDswjRic7b68zXuVpaVzAKQKx5UgJqUxCl
46DB2y5vzA44fx+Pz7e/UIEHlqo9i7MzLfy6t75kYdY0/wxIn8hLFSOjLjvLaydr4W1YtlR2moSJ
lThHQ2416fMl/1DZ5bjkXq4eT+PXM9fQg4QgnV2TEyiq5o5Zm4Sef5DUk+3Ym7np0MStPg30HBQL
w8ZaOvIy53I5MsGxCCJ8bvcauDS7QaNtVb7DLU+VmVCFWAt/oxtvHWYXis8ZWQHzkofEqPHcHYR/
yF67WsTl4ZSdysU9BsiiapGkU2uZFFwrUZuOureraOXu/NjtCLtx883CZ3ZMKN89+PQVWkQD0TgH
e7jpzxyOHFkNG7bztA4Lwbucx/MggOFJKg2C1k/EMjYm/0ZJN97ggqWfwnLJJMMxrFMWxnhECmi3
CdbKR7Z8Tr4IjrVnT/CIwmAsyI6EifwdNk3PyRxYhBDaM2ECWJCFHmK6zlXwceI28K4SsYtKPkjz
nse3P4mmjbYlJnUcEfGgnICgt61RQrkiUWh1LbMleQBy3NJPTeVc/CsU2+sP7/RYrW+ykU3qqwEY
JBUusx1v9WoCiRrFbQF74f2gdcfBx6xjszEjP3UeBbVxnSxZ3dhKxap2HEX0lqayeRhQ2leMKVFS
W/NOUGxo7dRnjLnxL9VgRk1ulVhREAbtn+Ro3kmo7iDMIl8I88BAe6Eq3b4xilB/IMCuAPE+jHM5
SXWhL396Uf1YT0hGG4oQ4B2oZK4aCZ3x09vSeVZqBlPYfNeTg9XLGIIMlh8HnMKgrpEcfiV6fu/G
ixl+KwWpo6dgLs4xvP5RqV82xm55TDfOEfuJxAdtc8gFYU2v6gEX1hWqp7Oq6pdX+V3H+m23z39f
iGnt8DTLqD71fx89bKLigarAHcd7HX02//RIGt6HQU03CHk+3EiKqgKBLR7utDM8205mqlRYmDgW
XItIttke7ZXhvXPlZ072+0UXj5AOV96Kmq4l6DE436a6iKlnbpSCSKf5MQ2zUdKD542nH4/18sHy
SBKHT/V8NJioXiTBTzoXXd1OVg9mS1aYsJznLQltk3erxtS8Kr/nSYN8jqwOCjf+NDjese+HdoVd
il5Y8Jg4FwDoJj/RVBiB3YBM496fr10SiuEbWDJ3ADfERf+YRMEHyTUrl4DbZtm2xNzoBBbdJAQ+
0cPJIKplxVOSp4jS5U35qHbUw2PZ15FPqc9zuBzTVjwYt2MyVSE0M0g2tqVEkqrx/XLGepNdDeKD
4jQ7O1b/YF648jL/cKJO6tXqfoXIPwRTGRChnu0WDhP8N4txP9wq9uD9lR9zl3XX+I3LgGUOZX3+
Y4tIsy3dun++Mm6gIJpf/WukKvSmvpUSxMg6lrpC6cwlY62HWMMUN8t/gV1GnaDLu3UApWsIMc/v
6nPx/jcdpGXa0N9hPY6jbIIoNnrZCAEgKFAVHaGQDrZrY3lZUROtyQyqyfvlUN0Ck0IqfnD1dcGB
bAXhadqO9ejObZysLNJ5vfOB77AeNu0zmB7F6aiuHQD7uhxrPPdFZhJSHmcBGs51QC93LsY9+/u+
0luJL//hJRlYrvYt4u9mNWBv7BV7HXMM51sgGMbpSQPuzSKPktJ9x4W1mR0rDaF6ENa0bGP1O/zr
eFJOIItOVpNrO3ksKouZXMwF+9qhFZua3h+SsScMN79Fs5+0hw72iIm2PHLTBDzDeXXGl3sUMx5W
wcnDr5dWSbAI/DtKsREbDgwKdBEJyQ1CK+4a0IRCyVeZkAIZ/gL6YiSwwXMkMf3n6lpCGWgnIyAr
y6yM5mpdxtsxNgurIz4aTi7dco8zdy0DhoWtAyVoUdODaD/imTQe00GpJTMMnnRkkr8TlilIMFUc
lqt9rkfduYgDy+wenqfcxD3CvgsOHvrjm4hsiIAI0jBqmSe6paPwH2WNULkNIN9MX3DAT6HocUfk
FSTtj2JcHQT6K0x/hh2t5h6ALBku4LaJAejjUTe9keeg+KuAurfTbW6FSEkiRVx4nW3ETfT6UG8q
amvnqI7BCIl2w2AVk24ZVxE1h0Yws2bko+85BHbKLwxvFiNDa3fzfFJKsVfRglgT7fXca6PMC/bx
gBa8NAR/tYzZGyU3fOS1ed03WytjbEiJjMmo7cJWEkpaIivT1OwmLXgwEU02C/UsoPdX9pFN/Aoj
dUA/kIeRzyll5b/wtZD6dxvcA7DBFPwNxHNkMydEkwxVx2dzRfx4n3DKGDLMXKKcqq3dzMKYakJt
CBZRWynitGg68aoQ8iFKOXuXLsPpIVJ+HPMkq76ykdlP2fQYTdl+xXzpiKusSMGLeXw1L0b1TfsA
ReyQ/dfsH4fFh24/aD/Onmmt1rbLpWRHrt87uNcKaZjmHIPZLkND5bsyIYctxUpxBdDJrYggo6ne
bHsxxR0/iY4rlGhaVz9mcJA9INC4pcx/C129h+XfN6/QiMtQg+h+x3LuXJS7e70eE+wXsVrY91R6
2iISnY/HGskfAWugOWqj5KmLZEcnQyZpf/fnN4PZajTqoJ7L/n20FQYnQmrZBgtyxyt+8ZTECSAq
sgeer7U69CA2yI3kkgmksK9fUzQGDGAtNcuJ2svgAreEfjRg/jYLtC9euF9OQlh2TS2DJiwPe8im
En7lEZtZskYAnE4ZdjyExhzvl53uQRpbyganmmaubmGv1JcAKA2FXcHNDzqf2s8qsz4OD4GwEhBA
pSH0I/2KfGHjqof3SqVDPOTOcJmoDHl0V6Uw9YGGKsSeaGZ3c3tNUG49dAJOCctYA2gBcXsaNNyd
uKPJ00mN0/W4ffgjUfFUTYsSVUF1qnoieaWRVAAQGM2pyD5iO88xN6UrSi/lsR756oa3pAmxzLeM
YP/kFge29vKeTh168KSS95mYRDhsLj/GjG5pWmb9ZnbEiZ+wVAi5f3Ba1cT9W6buXUUwXYRSyopB
KheF2qwSrw6WT1EFfx86UsdPdzYxi5a/ABLDHc+0BbTHn4f2mlotytp8nIN8BK/5PeyxOLh2bSvN
O5yqSqOjO7eQLEAn+kT1JwusapjXr8/AZG0O1ahzy7JEuIAr3RFok0lu6JVtnDIYQn5y+Pgg5bQ6
d16VhsGvJrepTFOlO4bcK5rmVIWj4nBIA1cHH/30LJJX4kBFjguQRKKub4I6aqibWSgGdTe4nW1P
2DdXjByhOdd+aMhDUTemYq6kFcGy2hNY2lG6y+QobBMyX+u3ttE+hcyptoH485JVjFQedkrL9meG
oOOhW2WmbBLUfDdCx3p0j2JadnRs+SJYlCkV1aJ8vSZPDO31epI90JfnZH9DUGmZm1KyZOanOl2U
sGthbR9x3stRUUfV2Ec4AnYq0yrZSQM7PL8FJ3dhj3WQqHecGC0JUmuW41g0yD17ha2ZZsiO2Rd5
DtGu0couJCx2jBC6/AV2oSI3Moy2ez73JCb4iVrNf4mX
`protect end_protected
